* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__oai33_1.ext - technology: gf180mcuD

.option scale=5n

X0 a_n200_690# B a_n370_690# VDD pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X1 a_n370_180# C OUT VSS nfet_03v3 ad=9.35n pd=0.28m as=17n ps=0.54m w=170 l=60
X2 a_n370_180# E VSS VSS nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X3 a_n370_690# C OUT VDD pfet_03v3 ad=18.7n pd=0.45m as=34n ps=0.88m w=340 l=60
X4 a_310_690# E a_140_690# VDD pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X5 VSS D a_n370_180# VSS nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X6 VSS F a_n370_180# VSS nfet_03v3 ad=17n pd=0.54m as=9.35n ps=0.28m w=170 l=60
X7 OUT F a_310_690# VDD pfet_03v3 ad=34n pd=0.88m as=18.7n ps=0.45m w=340 l=60
X8 a_n370_180# A OUT VSS nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X9 a_140_690# D VDD VDD pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X10 VDD A a_n200_690# VDD pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X11 OUT B a_n370_180# VSS nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
C0 F VDD 0.09613f
C1 A VDD 0.1093f
C2 C A 0.02542f
C3 a_310_690# F 0
C4 C VDD 0.11379f
C5 a_310_690# VDD 0.01042f
C6 D OUT 0.04618f
C7 D B 0.02346f
C8 a_n370_180# OUT 0.27551f
C9 D E 0.06224f
C10 B a_n370_180# 0.01381f
C11 a_n200_690# VDD 0.011f
C12 E a_n370_180# 0.04792f
C13 a_140_690# OUT 0.01568f
C14 F OUT 0.05506f
C15 E F 0.06521f
C16 A OUT 0.0953f
C17 a_n370_690# VDD 0.01042f
C18 B A 0.06224f
C19 C a_n370_690# 0.0028f
C20 OUT VDD 0.36514f
C21 C OUT 0.22193f
C22 A E 0.02346f
C23 B VDD 0.09001f
C24 C B 0.07167f
C25 D a_n370_180# 0.12372f
C26 E VDD 0.10378f
C27 a_310_690# OUT 0.01597f
C28 a_310_690# E 0.00187f
C29 D a_140_690# 0.00156f
C30 D F 0.02542f
C31 a_n200_690# OUT 0.01568f
C32 B a_n200_690# 0.00156f
C33 a_n370_180# F 0.00529f
C34 D A 0.06224f
C35 D VDD 0.09371f
C36 A a_n370_180# 0.03452f
C37 a_n370_180# VDD 0.0041f
C38 C a_n370_180# 0.00483f
C39 a_n370_690# OUT 0.01597f
C40 B OUT 0.18496f
C41 a_140_690# VDD 0.011f
C42 E OUT 0.12283f
C43 OUT VSS 0.52966f
C44 F VSS 0.37682f
C45 E VSS 0.27402f
C46 D VSS 0.29097f
C47 A VSS 0.26783f
C48 B VSS 0.28758f
C49 C VSS 0.33492f
C50 VDD VSS 2.76557f
C51 a_n370_180# VSS 0.76901f **FLOATING
