* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.2.ext - technology: gf180mcuC

X0 a_1160_210# C1.t0 OUT.t1 VDD.t5 pfet_03v3 ad=0.85p pd=4.4u as=0.595p ps=2.4u w=1.7u l=0.3u
X1 X2.t1 a_250_210# a_590_210# VSS.t9 nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 X0.t1 a_250_210# a_1160_210# VSS.t8 nfet_03v3 ad=0.5525p pd=3u as=0.32p ps=1.65u w=0.85u l=0.3u
X3 X2.t0 C0.t0 a_590_210# VDD.t2 pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
X4 a_n90_210# C1.t1 VSS.t3 VSS.t2 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 X0.t0 C0.t1 a_1160_210# VDD.t7 pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
X6 a_250_210# C0.t2 VSS.t5 VSS.t4 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 OUT.t0 C1.t2 a_590_210# VSS.t1 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 a_n90_210# C1.t3 VDD.t4 VDD.t3 pfet_03v3 ad=1.02p pd=4.6u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_250_210# C0.t3 VDD.t1 VDD.t0 pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X10 OUT.t2 a_n90_210# a_590_210# VDD.t6 pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X11 a_590_210# C0.t4 X3.t0 VSS.t7 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# C0.t5 X1.t0 VSS.t0 nfet_03v3 ad=0.32p pd=1.65u as=0.425p ps=2.7u w=0.85u l=0.3u
X13 a_590_210# a_250_210# X3.t1 VDD.t9 pfet_03v3 ad=0.595p pd=2.4u as=0.87p ps=4.5u w=1.7u l=0.3u
X14 a_1160_210# a_n90_210# OUT.t3 VSS.t6 nfet_03v3 ad=0.6025p pd=3.2u as=0.2975p ps=1.55u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# X1.t1 VDD.t8 pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
C0 X3 a_250_210# 0.38226f
C1 a_n90_210# OUT 0.1469f
C2 X2 C0 0.12331f
C3 VDD X1 0.05854f
C4 X3 X2 0.01084f
C5 X0 X1 0.01101f
C6 a_1160_210# a_250_210# 0.02157f
C7 a_590_210# a_250_210# 0.03134f
C8 C0 OUT 0.00857f
C9 X1 C1 0.0177f
C10 C0 a_n90_210# 0.52899f
C11 VDD a_250_210# 0.90117f
C12 X3 OUT 0
C13 a_1160_210# X2 0.00111f
C14 a_590_210# X2 0.24495f
C15 X3 a_n90_210# 0.01988f
C16 X0 a_250_210# 0.00583f
C17 VDD X2 0.06725f
C18 a_250_210# C1 0.03025f
C19 a_1160_210# OUT 0.22347f
C20 a_590_210# OUT 0.34464f
C21 a_1160_210# a_n90_210# 0.14865f
C22 X3 C0 0.05504f
C23 a_590_210# a_n90_210# 0.10406f
C24 X2 C1 0.01941f
C25 VDD OUT 0.05981f
C26 VDD a_n90_210# 0.51229f
C27 X0 OUT 0.00308f
C28 X0 a_n90_210# 0.05776f
C29 a_1160_210# C0 0.16894f
C30 a_590_210# C0 0.24844f
C31 OUT C1 0.08109f
C32 a_n90_210# C1 1.09594f
C33 VDD C0 0.41598f
C34 X3 a_1160_210# 0
C35 X3 a_590_210# 0.33193f
C36 X1 a_250_210# 0.03933f
C37 X0 C0 0.08388f
C38 X3 VDD 0.06719f
C39 X2 X1 0.37477f
C40 C0 C1 0.05297f
C41 a_1160_210# a_590_210# 0.03595f
C42 X3 C1 0.01791f
C43 a_1160_210# VDD 0.11343f
C44 VDD a_590_210# 0.28685f
C45 X1 OUT 0
C46 X1 a_n90_210# 0.01895f
C47 X2 a_250_210# 0.03826f
C48 a_1160_210# X0 0.20157f
C49 X0 a_590_210# 0.39419f
C50 a_1160_210# C1 0.55003f
C51 a_590_210# C1 0.05053f
C52 X0 VDD 0.06734f
C53 VDD C1 0.54837f
C54 X1 C0 0.05434f
C55 a_250_210# OUT 0
C56 a_250_210# a_n90_210# 0.08779f
C57 X0 C1 0.0258f
C58 X2 OUT 0
C59 X2 a_n90_210# 0.01989f
C60 a_250_210# C0 0.3665f
C61 a_1160_210# X1 0.33285f
C62 a_590_210# X1 0.05209f
R0 C1.n0 C1.t2 90.406
R1 C1 C1.n0 71.1138
R2 C1.n1 C1.t1 36.5005
R3 C1.n0 C1.t0 34.6755
R4 C1.n1 C1.t3 29.8088
R5 C1 C1.n1 12.5005
R6 OUT.n2 OUT.n1 6.8405
R7 OUT.n3 OUT.n2 4.5005
R8 OUT.n1 OUT.t3 3.1505
R9 OUT.n2 OUT.n0 2.21083
R10 OUT.n1 OUT.t0 2.03874
R11 OUT.n0 OUT.t1 1.7505
R12 OUT.n0 OUT.t2 1.13285
R13 OUT OUT.n3 0.03425
R14 OUT.n3 OUT 0.03425
R15 VDD.t8 VDD.t2 578.125
R16 VDD.t7 VDD.n2 570.312
R17 VDD.t3 VDD.n7 398.438
R18 VDD.t6 VDD.t5 312.5
R19 VDD.t2 VDD.t9 312.5
R20 VDD.n3 VDD.t8 304.688
R21 VDD.n6 VDD.t9 273.438
R22 VDD.t0 VDD.n6 257.812
R23 VDD.t5 VDD.n1 176.863
R24 VDD.n7 VDD.t0 132.812
R25 VDD VDD.t3 98.538
R26 VDD.n2 VDD.n1 12.6005
R27 VDD.n4 VDD.n3 12.6005
R28 VDD.n6 VDD.n5 12.6005
R29 VDD.n7 VDD.n0 12.6005
R30 VDD.n2 VDD.t6 7.813
R31 VDD.n3 VDD.t7 7.813
R32 VDD VDD.t4 3.3014
R33 VDD.n0 VDD.t1 3.29819
R34 VDD.n5 VDD.n4 0.604786
R35 VDD.n4 VDD.n1 0.238357
R36 VDD VDD.n0 0.199786
R37 VDD.n5 VDD.n0 0.161214
R38 X2.n0 X2.t1 10.4272
R39 X2.n1 X2.n0 4.57
R40 X2.n0 X2.t0 4.351
R41 X2 X2.n1 0.0275
R42 X2.n1 X2 0.0275
R43 VSS.t9 VSS.t0 1908.73
R44 VSS.n2 VSS.t1 1367.06
R45 VSS.n7 VSS.t7 1109.13
R46 VSS.t2 VSS.n8 1057.54
R47 VSS.t1 VSS.t6 1031.75
R48 VSS.t0 VSS.t8 1031.75
R49 VSS.n3 VSS.t9 748.016
R50 VSS.n8 VSS.t4 696.429
R51 VSS.t4 VSS.n7 644.841
R52 VSS.t6 VSS.n1 604.028
R53 VSS.t8 VSS.n2 541.668
R54 VSS VSS.t2 448.892
R55 VSS.n3 VSS.t7 283.731
R56 VSS.n2 VSS.n1 10.4005
R57 VSS.n4 VSS.n3 10.4005
R58 VSS.n7 VSS.n6 10.4005
R59 VSS.n8 VSS.n0 10.4005
R60 VSS.n5 VSS.t5 8.61774
R61 VSS VSS.t3 8.61774
R62 VSS.n4 VSS.n1 0.527643
R63 VSS VSS.n0 0.186929
R64 VSS.n6 VSS.n4 0.174071
R65 VSS.n6 VSS.n5 0.1355
R66 VSS.n5 VSS.n0 0.0326429
R67 X0.n0 X0.t1 10.4272
R68 X0.n1 X0.n0 4.57
R69 X0.n0 X0.t0 4.351
R70 X0 X0.n1 0.0275
R71 X0.n1 X0 0.0275
R72 C0.n1 C0.t4 45.6255
R73 C0.n0 C0.t5 45.6255
R74 C0.n3 C0.t2 36.777
R75 C0.n1 C0.t0 30.4172
R76 C0.n0 C0.t1 30.4172
R77 C0.n3 C0.t3 30.0854
R78 C0.n2 C0.n0 13.3212
R79 C0.n4 C0.n3 12.5005
R80 C0.n2 C0.n1 12.5005
R81 C0.n4 C0.n2 0.808357
R82 C0 C0.n4 0.03425
R83 X3.n0 X3.t0 9.31403
R84 X3.n1 X3.n0 4.5685
R85 X3.n0 X3.t1 3.73335
R86 X3 X3.n1 0.0275
R87 X3.n1 X3 0.0275
R88 X1.n0 X1.t0 9.31403
R89 X1.n1 X1.n0 4.5685
R90 X1.n0 X1.t1 3.73335
R91 X1 X1.n1 0.0275
R92 X1.n1 X1 0.0275
C63 OUT VSS 0.12063f
C64 X0 VSS 0.11279f
C65 X1 VSS 0.09904f
C66 X2 VSS 0.10766f
C67 X3 VSS 0.12007f
C68 C0 VSS 1.05023f
C69 C1 VSS 1.39324f
C70 VDD VSS 5.51923f
C71 a_1160_210# VSS 0.71666f **FLOATING
C72 a_590_210# VSS 0.36135f **FLOATING
C73 a_n90_210# VSS 1.23339f **FLOATING
C74 a_250_210# VSS 1.3406f **FLOATING
