* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__oai33_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__oai33_1 A B C D E F OUT VDD VSS
X0 a_n200_690# B a_n370_690# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 a_n370_180# C OUT VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X2 a_n370_180# E VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 a_n370_690# C OUT VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 a_310_690# E a_140_690# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 VSS D a_n370_180# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X6 VSS F a_n370_180# VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X7 OUT F a_310_690# VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X8 a_n370_180# A OUT VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X9 a_140_690# D VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X10 VDD A a_n200_690# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X11 OUT B a_n370_180# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
C0 a_140_690# VDD 0.011f
C1 OUT D 0.04618f
C2 A C 0.02542f
C3 a_310_690# F 0
C4 A D 0.06224f
C5 E a_n370_180# 0.04792f
C6 VDD a_n370_690# 0.01042f
C7 B a_n370_180# 0.01381f
C8 E F 0.06521f
C9 VDD a_n370_180# 0.0041f
C10 A OUT 0.0953f
C11 D E 0.06224f
C12 OUT a_310_690# 0.01597f
C13 C B 0.07167f
C14 VDD F 0.09613f
C15 B D 0.02346f
C16 VDD C 0.11379f
C17 VDD D 0.09371f
C18 OUT a_n200_690# 0.01568f
C19 OUT E 0.12283f
C20 a_140_690# D 0.00156f
C21 OUT B 0.18496f
C22 A E 0.02346f
C23 C a_n370_690# 0.0028f
C24 OUT VDD 0.36514f
C25 a_310_690# E 0.00187f
C26 A B 0.06224f
C27 a_140_690# OUT 0.01568f
C28 A VDD 0.1093f
C29 a_n370_180# F 0.00529f
C30 C a_n370_180# 0.00483f
C31 VDD a_310_690# 0.01042f
C32 D a_n370_180# 0.12372f
C33 B a_n200_690# 0.00156f
C34 OUT a_n370_690# 0.01597f
C35 VDD a_n200_690# 0.011f
C36 D F 0.02542f
C37 VDD E 0.10378f
C38 OUT a_n370_180# 0.27551f
C39 VDD B 0.09001f
C40 A a_n370_180# 0.03452f
C41 OUT F 0.05506f
C42 OUT C 0.22193f
C43 OUT VSS 0.52966f
C44 F VSS 0.37682f
C45 E VSS 0.27402f
C46 D VSS 0.29097f
C47 A VSS 0.26783f
C48 B VSS 0.28758f
C49 C VSS 0.33492f
C50 VDD VSS 2.76557f
C51 a_n370_180# VSS 0.76901f
.ends gf180mcu_osu_sc_gp9t3v3__oai33_1

