* OAI33 functional verification (LVS-extracted netlist, no parasitics)
* Logic: Y = ~((A|B|C) & (D|E|F))

************** MODELS **************
.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

************** SUBCKT **************
* Pin order: VDD A B C D E F OUT VSS
.subckt gf180mcu_osu_sc_gp9t3v3__oai33_1 VDD A B C D E F OUT VSS

X0  a_n200_690#  B  a_n370_690#  VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1  a_n370_180#  C  OUT         VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p  ps=2.7u  w=0.85u l=0.3u
X2  a_n370_180#  E  VSS         VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3  a_n370_690#  C  OUT         VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p   ps=4.4u w=1.7u l=0.3u
X4  a_310_690#   E  a_140_690#  VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5  VSS          D  a_n370_180# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X6  VSS          F  a_n370_180# VSS nfet_03v3 ad=0.425p  pd=2.7u  as=0.23375p ps=1.4u w=0.85u l=0.3u
X7  OUT          F  a_310_690#  VDD pfet_03v3 ad=0.85p   pd=4.4u  as=0.4675p ps=2.25u w=1.7u l=0.3u
X8  a_n370_180#  A  OUT         VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X9  a_140_690#   D  VDD         VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X10 VDD          A  a_n200_690# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X11 OUT          B  a_n370_180# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u

.ends gf180mcu_osu_sc_gp9t3v3__oai33_1

************** PARAMS **************
.param VDDval = 3.3
.param trise  = 500p
.param tfall  = 500p
.param tpulse = 50n     
.param tdelay = 0

************** SOURCES **************
VDD   VDD  0  {VDDval}

* Input stimuli pakai counter style
* Period tiap input = 2x dari input sebelumnya
VA  A  0  PULSE(0 {VDDval} {tdelay} {trise} {tfall} {8*tpulse} {16*tpulse})
VB  B  0  PULSE(0 {VDDval} {tdelay} {trise} {tfall} {4*tpulse} {8*tpulse})
VC  C  0  PULSE(0 {VDDval} {tdelay} {trise} {tfall} {2*tpulse} {4*tpulse})
VD  D  0  PULSE(0 {VDDval} {tdelay} {trise} {tfall} {1*tpulse} {2*tpulse})
VE  E  0  PULSE(0 {VDDval} {tdelay} {trise} {tfall} {0.5*tpulse} {1*tpulse})
VF  F  0  PULSE(0 {VDDval} {tdelay} {trise} {tfall} {0.25*tpulse} {0.5*tpulse})

* DUT
XU1 VDD A B C D E F OUT 0 gf180mcu_osu_sc_gp9t3v3__oai33_1


.control
    run
    set color0=white
    set color1=black
    set xbrushwidth=3
    tran 0.01ns 810ns
    plot out a+4 b+8 c+12 d+16 e+20 f+24
.endc