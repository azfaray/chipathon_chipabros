* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__oai33_1.2.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__oai33_1 A B C D E F OUT VDD VSS

X0 a_n200_690# B.t0 a_n370_690# VDD.t7 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 a_n370_180# C.t0 OUT.t1 VSS.t2 nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X2 a_n370_180# E.t0 VSS.t1 VSS.t0 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 a_n370_690# C.t1 OUT.t0 VDD.t3 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 a_310_690# E.t1 a_140_690# VDD.t2 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 VSS.t4 D.t0 a_n370_180# VSS.t3 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X6 VSS.t6 F.t0 a_n370_180# VSS.t5 nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X7 OUT.t2 F.t1 a_310_690# VDD.t4 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X8 a_n370_180# A.t0 OUT.t3 VSS.t7 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X9 a_140_690# D.t1 VDD.t1 VDD.t0 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X10 VDD.t6 A.t1 a_n200_690# VDD.t5 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X11 OUT.t4 B.t1 a_n370_180# VSS.t8 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
C0 E a_310_690# 0.00187f
C1 VDD a_n370_180# 0.0041f
C2 VDD D 0.09371f
C3 E F 0.06521f
C4 C a_n370_690# 0.0028f
C5 a_n370_180# D 0.12372f
C6 VDD OUT 0.36514f
C7 VDD a_n200_690# 0.011f
C8 F a_310_690# 0
C9 VDD A 0.1093f
C10 a_n370_180# OUT 0.27551f
C11 a_n370_180# A 0.03452f
C12 D OUT 0.04618f
C13 VDD B 0.09001f
C14 D A 0.06224f
C15 VDD E 0.10378f
C16 a_n370_180# B 0.01381f
C17 OUT a_n200_690# 0.01568f
C18 a_n370_180# E 0.04792f
C19 A OUT 0.0953f
C20 VDD C 0.11379f
C21 B D 0.02346f
C22 VDD a_310_690# 0.01042f
C23 E D 0.06224f
C24 C a_n370_180# 0.00483f
C25 VDD a_n370_690# 0.01042f
C26 B OUT 0.18496f
C27 B a_n200_690# 0.00156f
C28 VDD F 0.09613f
C29 E OUT 0.12283f
C30 B A 0.06224f
C31 VDD a_140_690# 0.011f
C32 a_n370_180# F 0.00529f
C33 E A 0.02346f
C34 C OUT 0.22193f
C35 OUT a_310_690# 0.01597f
C36 D F 0.02542f
C37 C A 0.02542f
C38 D a_140_690# 0.00156f
C39 OUT a_n370_690# 0.01597f
C40 F OUT 0.05506f
C41 C B 0.07167f
C42 OUT a_140_690# 0.01568f
R0 B.n0 B.t0 46.2338
R1 B.n0 B.t1 21.2922
R2 B.n1 B.n0 12.5005
R3 B B.n1 0.0275
R4 B.n1 B 0.0275
R5 VDD.t2 VDD.t0 265.625
R6 VDD.t5 VDD.n5 226.562
R7 VDD.t7 VDD.n6 164.062
R8 VDD.n7 VDD.t7 164.062
R9 VDD.n6 VDD.t5 101.562
R10 VDD.n7 VDD.t3 101.562
R11 VDD.n1 VDD.t4 67.6105
R12 VDD.n5 VDD.t0 39.063
R13 VDD.n1 VDD.t2 32.0719
R14 VDD.n5 VDD.n4 12.6005
R15 VDD.n6 VDD.n0 12.6005
R16 VDD VDD.n7 12.6005
R17 VDD.n4 VDD.n1 3.65344
R18 VDD.n3 VDD.n2 2.9425
R19 VDD.n2 VDD.t1 1.13285
R20 VDD.n2 VDD.t6 1.13285
R21 VDD VDD.n0 0.1355
R22 VDD.n3 VDD.n0 0.0969286
R23 VDD.n4 VDD.n3 0.0390714
R24 C.n0 C.t0 36.5005
R25 C.n0 C.t1 29.8088
R26 C.n1 C.n0 12.5005
R27 C C.n1 0.0275
R28 C.n1 C 0.0275
R29 OUT.n1 OUT.t1 8.45574
R30 OUT.n1 OUT.n0 6.9575
R31 OUT.n4 OUT.n3 4.7075
R32 OUT.n3 OUT.t2 3.08219
R33 OUT.n2 OUT.t0 3.08219
R34 OUT.n0 OUT.t3 2.03874
R35 OUT.n0 OUT.t4 2.03874
R36 OUT.n3 OUT.n2 1.8365
R37 OUT.n2 OUT.n1 0.5585
R38 OUT OUT.n4 0.03425
R39 OUT.n4 OUT 0.03425
R40 VSS.t0 VSS.t3 876.985
R41 VSS.n3 VSS.t5 799.604
R42 VSS.t7 VSS.n7 748.016
R43 VSS.t8 VSS.n8 541.668
R44 VSS.n9 VSS.t8 541.668
R45 VSS.n8 VSS.t7 335.317
R46 VSS.n9 VSS.t2 335.317
R47 VSS.t5 VSS.n2 294.13
R48 VSS.n7 VSS.t3 128.969
R49 VSS.n3 VSS.t0 77.3815
R50 VSS.n4 VSS.n3 10.4005
R51 VSS.n7 VSS.n6 10.4005
R52 VSS.n8 VSS.n0 10.4005
R53 VSS VSS.n9 10.4005
R54 VSS.n2 VSS.t6 8.63702
R55 VSS.n5 VSS.n1 6.5165
R56 VSS.n1 VSS.t1 2.03874
R57 VSS.n1 VSS.t4 2.03874
R58 VSS.n4 VSS.n2 0.1355
R59 VSS.n6 VSS.n0 0.1355
R60 VSS VSS.n0 0.1355
R61 VSS.n6 VSS.n5 0.0712143
R62 VSS.n5 VSS.n4 0.0647857
R63 E.n0 E.t0 37.1088
R64 E.n0 E.t1 30.4172
R65 E.n1 E.n0 12.5005
R66 E E.n1 0.0275
R67 E.n1 E 0.0275
R68 D.n0 D.t1 46.2338
R69 D.n0 D.t0 21.2922
R70 D.n1 D.n0 12.5005
R71 D D.n1 0.0275
R72 D.n1 D 0.0275
R73 F.n0 F.t1 46.2338
R74 F.n0 F.t0 21.2922
R75 F.n1 F.n0 12.5005
R76 F F.n1 0.0275
R77 F.n1 F 0.0275
R78 A.n0 A.t0 37.1088
R79 A.n0 A.t1 30.4172
R80 A.n1 A.n0 12.5005
R81 A A.n1 0.0275
R82 A.n1 A 0.0275
C43 OUT VSS 0.52966f
C44 F VSS 0.37682f
C45 E VSS 0.27402f
C46 D VSS 0.29097f
C47 A VSS 0.26783f
C48 B VSS 0.28758f
C49 C VSS 0.33492f
C50 VDD VSS 2.76557f
C51 a_n370_180# VSS 0.76901f
.ends gf180mcu_osu_sc_gp9t3v3__oai33_1