* NGSPICE file created from MUX4.ext - technology: gf180mcuC

.subckt MUX4 OUT X0 X1 X3 X2 C1 C0 VDD VSS
X0 a_1160_210# C1 OUT VDD pfet_03v3 ad=0.85p pd=4.4u as=0.595p ps=2.4u w=1.7u l=0.3u
X1 X2 a_250_210# a_590_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 X0 a_250_210# a_1160_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.32p ps=1.65u w=0.85u l=0.3u
X3 X2 C0 a_590_210# VDD pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X4 a_n90_210# C1 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 X0 C0 a_1160_210# VDD pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X6 a_250_210# C0 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 OUT C1 a_590_210# VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 a_n90_210# C1 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_250_210# C0 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X10 OUT a_n90_210# a_590_210# VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X11 a_590_210# C0 X3 VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# C0 X1 VSS nfet_03v3 ad=0.32p pd=1.65u as=0.425p ps=2.7u w=0.85u l=0.3u
X13 a_590_210# a_250_210# X3 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X14 a_1160_210# a_n90_210# OUT VSS nfet_03v3 ad=0.6025p pd=3.2u as=0.2975p ps=1.55u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# X1 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
C0 OUT a_590_210# 0.34464f
C1 X3 VDD 0.09082f
C2 X2 a_590_210# 0.22961f
C3 a_1160_210# a_590_210# 0.03595f
C4 a_250_210# VDD 0.90082f
C5 a_n90_210# OUT 0.1469f
C6 X2 a_n90_210# 0.02067f
C7 a_1160_210# a_n90_210# 0.14845f
C8 X1 a_250_210# 0.04064f
C9 OUT C1 0.07582f
C10 C0 X0 0.08405f
C11 X2 C1 0.01928f
C12 a_1160_210# C1 0.53587f
C13 X0 a_590_210# 0.37242f
C14 a_n90_210# X0 0.05962f
C15 C0 VDD 0.41628f
C16 X2 OUT 0
C17 a_1160_210# OUT 0.22347f
C18 VDD a_590_210# 0.28422f
C19 a_1160_210# X2 0.00111f
C20 a_250_210# X3 0.37991f
C21 a_n90_210# VDD 0.51226f
C22 X0 C1 0.02056f
C23 X1 C0 0.06472f
C24 X1 a_590_210# 0.03496f
C25 VDD C1 0.42961f
C26 OUT X0 0.00299f
C27 X1 a_n90_210# 0.01914f
C28 a_1160_210# X0 0.20363f
C29 C0 X3 0.04882f
C30 OUT VDD 0.05981f
C31 X3 a_590_210# 0.35452f
C32 a_250_210# C0 0.3665f
C33 X2 VDD 0.06601f
C34 a_1160_210# VDD 0.11048f
C35 a_250_210# a_590_210# 0.03014f
C36 X1 C1 0.01724f
C37 a_n90_210# X3 0.01961f
C38 a_n90_210# a_250_210# 0.08868f
C39 X1 OUT 0
C40 X2 X1 0.37197f
C41 a_1160_210# X1 0.32933f
C42 X3 C1 0.01769f
C43 VDD X0 0.06464f
C44 a_250_210# C1 0.02985f
C45 C0 a_590_210# 0.25009f
C46 OUT X3 0
C47 X2 X3 0.0012f
C48 a_1160_210# X3 0
C49 a_250_210# OUT 0
C50 a_n90_210# C0 0.52899f
C51 X2 a_250_210# 0.03943f
C52 a_1160_210# a_250_210# 0.02157f
C53 X1 X0 0.01083f
C54 a_n90_210# a_590_210# 0.10428f
C55 X1 VDD 0.05717f
C56 C0 C1 0.05224f
C57 C1 a_590_210# 0.04739f
C58 a_250_210# X0 0.00583f
C59 a_n90_210# C1 1.09377f
C60 OUT C0 0.00857f
C61 X2 C0 0.1344f
C62 a_1160_210# C0 0.16894f
C63 OUT VSS 0.12063f
C64 X0 VSS 0.11727f
C65 X1 VSS 0.09987f
C66 X2 VSS 0.11206f
C67 X3 VSS 0.12356f
C68 C0 VSS 1.0511f
C69 C1 VSS 1.35886f
C70 VDD VSS 5.40677f
C71 a_1160_210# VSS 0.72049f
C72 a_590_210# VSS 0.35695f
C73 a_n90_210# VSS 1.23402f
C74 a_250_210# VSS 1.33965f
.ends
