* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__aoi33_1.2.ext - technology: gf180mcuD

X0 a_1310_210# F.t0 VSS.t7 VSS.t6 nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 OUT.t0 D.t0 a_1480_210# VSS.t0 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X2 a_1480_210# E.t0 a_1310_210# VSS.t4 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 a_1310_720# F.t1 OUT.t4 VDD.t8 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 a_1310_720# D.t1 OUT.t1 VDD.t0 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 a_1820_210# A.t0 OUT.t3 VSS.t1 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X6 OUT.t2 E.t1 a_1310_720# VDD.t3 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X7 VSS.t3 C.t0 a_1990_210# VSS.t2 nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X8 a_1990_210# B.t0 a_1820_210# VSS.t5 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X9 VDD.t2 A.t1 a_1310_720# VDD.t1 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X10 VDD.t7 C.t1 a_1310_720# VDD.t6 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X11 a_1310_720# B.t1 VDD.t5 VDD.t4 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
C0 F C 0
C1 F A 0
C2 a_1820_210# OUT 0.00354f
C3 VDD OUT 0.16592f
C4 a_1310_720# OUT 0.62324f
C5 D OUT 0.18649f
C6 B VDD 0.09805f
C7 a_1310_720# B 0.02283f
C8 E F 0.07113f
C9 a_1480_210# D 0.00297f
C10 B OUT 0.09467f
C11 E a_1310_210# 0.00297f
C12 F VDD 0.13074f
C13 F D 0
C14 F a_1310_720# 0.00167f
C15 a_1990_210# OUT 0.00297f
C16 a_1480_210# OUT 0.00316f
C17 a_1990_210# B 0.00297f
C18 F OUT 0.11804f
C19 C VDD 0.10876f
C20 a_1820_210# A 0.00297f
C21 A VDD 0.09996f
C22 a_1310_720# C 0.00167f
C23 F B 0
C24 a_1310_720# A 0.01969f
C25 D A 0.06819f
C26 a_1310_210# OUT 0.00232f
C27 E VDD 0.08723f
C28 E a_1310_720# 0.01759f
C29 E D 0.13834f
C30 C OUT 0.10022f
C31 A OUT 0.1684f
C32 C B 0.13834f
C33 A B 0.13834f
C34 a_1310_720# VDD 0.72085f
C35 D VDD 0.08675f
C36 E OUT 0.05861f
C37 a_1310_720# D 0.0172f
R0 F.n1 F.t0 35.7401
R1 F.n1 F.t1 29.0484
R2 F.n2 F.n1 8.0005
R3 F F.n2 4.5185
R4 F.n2 F.n0 0.0185
R5 VSS.t5 VSS.t1 876.985
R6 VSS.t6 VSS.t4 876.985
R7 VSS.n3 VSS.t2 748.016
R8 VSS.t0 VSS.n6 644.841
R9 VSS.n7 VSS.t0 593.255
R10 VSS.t2 VSS.n2 500.486
R11 VSS.t4 VSS.n7 283.731
R12 VSS.n6 VSS.t1 232.143
R13 VSS.n3 VSS.t5 128.969
R14 VSS.n8 VSS.t6 82.5815
R15 VSS.n4 VSS.n3 10.4005
R16 VSS.n6 VSS.n5 10.4005
R17 VSS.n7 VSS.n0 10.4005
R18 VSS VSS.t7 8.65952
R19 VSS.n2 VSS.t3 8.61774
R20 VSS.n9 VSS.n8 5.2005
R21 VSS.n8 VSS.n1 0.389389
R22 VSS.n5 VSS.n4 0.154786
R23 VSS.n5 VSS.n0 0.154786
R24 VSS.n9 VSS.n0 0.154786
R25 VSS.n4 VSS.n2 0.148357
R26 VSS VSS.n9 0.00371429
R27 D.n1 D.t1 45.6255
R28 D.n1 D.t0 20.6838
R29 D.n2 D.n1 8.0005
R30 D D.n2 4.51175
R31 D.n2 D.n0 0.0155
R32 OUT.n4 OUT.n1 6.8315
R33 OUT OUT.n5 4.523
R34 OUT.n3 OUT.t4 3.57419
R35 OUT.n3 OUT.n2 2.7085
R36 OUT.n1 OUT.t3 2.03874
R37 OUT.n1 OUT.t0 2.03874
R38 OUT.n2 OUT.t1 1.13285
R39 OUT.n2 OUT.t2 1.13285
R40 OUT.n5 OUT.n4 1.0565
R41 OUT.n4 OUT.n3 0.4505
R42 OUT.n5 OUT.n0 0.0305
R43 E.n1 E.t1 45.6255
R44 E.n1 E.t0 20.6838
R45 E.n2 E.n1 8.0005
R46 E E.n2 4.51175
R47 E.n2 E.n0 0.0155
R48 VDD.t4 VDD.t1 265.625
R49 VDD.t8 VDD.t3 265.625
R50 VDD.n4 VDD.t6 226.562
R51 VDD.t0 VDD.n8 195.312
R52 VDD.n9 VDD.t0 179.689
R53 VDD.t6 VDD.n3 161.044
R54 VDD.t3 VDD.n9 85.938
R55 VDD.n8 VDD.t1 70.313
R56 VDD.n4 VDD.t4 39.063
R57 VDD.n10 VDD.t8 29.738
R58 VDD.n5 VDD.n4 12.6005
R59 VDD.n8 VDD.n7 12.6005
R60 VDD.n9 VDD.n0 12.6005
R61 VDD VDD.n10 6.30371
R62 VDD.n3 VDD.t7 3.29819
R63 VDD.n6 VDD.n2 2.9425
R64 VDD.n2 VDD.t5 1.13285
R65 VDD.n2 VDD.t2 1.13285
R66 VDD.n10 VDD.n1 0.3505
R67 VDD.n7 VDD.n0 0.154786
R68 VDD VDD.n0 0.151571
R69 VDD.n5 VDD.n3 0.148357
R70 VDD.n7 VDD.n6 0.0840714
R71 VDD.n6 VDD.n5 0.0712143
R72 A.n1 A.t1 45.6255
R73 A.n1 A.t0 20.6838
R74 A.n2 A.n1 8.0005
R75 A A.n2 4.51175
R76 A.n2 A.n0 0.0155
R77 C.n1 C.t1 45.6255
R78 C.n1 C.t0 20.6838
R79 C.n2 C.n1 8.0005
R80 C C.n2 4.51175
R81 C.n2 C.n0 0.0155
R82 B.n0 B.t1 45.6255
R83 B.n0 B.t0 20.6838
R84 B.n1 B.n0 8.0005
R85 B B.n1 4.5005
C38 OUT VSS 0.42162f
C39 C VSS 0.3984f
C40 B VSS 0.30452f
C41 A VSS 0.30946f
C42 D VSS 0.30954f
C43 E VSS 0.32807f
C44 F VSS 0.39864f
C45 VDD VSS 2.84616f
C46 a_1990_210# VSS 0.00795f 
C47 a_1820_210# VSS 0.00738f 
C48 a_1480_210# VSS 0.00738f 
C49 a_1310_210# VSS 0.00795f 
C50 a_1310_720# VSS 0.07075f 
