VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__mux4_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__mux4_1 ;
  ORIGIN 1.700 0.000 ;
  SIZE 12.450 BY 6.350 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -1.700 3.150 10.750 6.350 ;
      LAYER Metal1 ;
        RECT -1.700 5.650 10.750 6.350 ;
        RECT -1.150 3.600 -0.900 5.650 ;
        RECT 0.550 3.600 0.800 5.650 ;
    END
  END VDD
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.350 3.350 10.650 3.850 ;
        RECT -1.050 2.950 -0.550 3.250 ;
      LAYER Metal2 ;
        RECT 10.300 3.400 10.700 3.800 ;
        RECT -1.000 3.250 -0.600 3.300 ;
        RECT -1.000 2.950 -0.550 3.250 ;
        RECT -1.000 1.900 -0.600 2.950 ;
        RECT 10.350 1.900 10.650 3.400 ;
        RECT -1.000 1.600 10.650 1.900 ;
    END
  END C1
  PIN C0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.295000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 2.850 1.100 3.350 ;
        RECT 3.600 2.850 3.900 3.350 ;
        RECT 6.450 2.850 6.750 3.350 ;
      LAYER Metal2 ;
        RECT 0.750 3.250 1.150 3.300 ;
        RECT 3.500 3.250 4.000 3.300 ;
        RECT 6.350 3.250 6.850 3.300 ;
        RECT 0.750 2.950 6.850 3.250 ;
        RECT 0.750 2.900 1.150 2.950 ;
        RECT 3.550 2.900 3.950 2.950 ;
        RECT 6.400 2.900 6.800 2.950 ;
    END
  END C0
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT -1.150 0.700 -0.900 1.900 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT -1.700 0.000 10.750 0.700 ;
    END
  END VSS
  PIN X0
    DIRECTION INPUT ;
    ANTENNADIFFAREA 1.672500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 4.000 7.350 5.300 ;
        RECT 7.000 3.700 7.500 4.000 ;
        RECT 7.100 1.050 7.350 3.700 ;
      LAYER Metal2 ;
        RECT 7.050 4.000 7.450 4.050 ;
        RECT 7.050 3.700 7.500 4.000 ;
        RECT 7.050 3.650 7.450 3.700 ;
    END
  END X0
  PIN X1
    DIRECTION INPUT ;
    ANTENNADIFFAREA 1.290000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 4.000 5.350 5.300 ;
        RECT 4.950 3.700 5.450 4.000 ;
        RECT 5.100 1.050 5.350 3.700 ;
      LAYER Metal2 ;
        RECT 5.000 4.000 5.400 4.050 ;
        RECT 5.000 3.700 5.450 4.000 ;
        RECT 5.000 3.650 5.400 3.700 ;
    END
  END X1
  PIN OUT
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.785000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.800 3.200 9.050 5.300 ;
        RECT 8.550 2.900 9.050 3.200 ;
        RECT 8.800 1.050 9.050 2.900 ;
      LAYER Metal2 ;
        RECT 8.600 2.850 9.050 3.250 ;
    END
  END OUT
  PIN X2
    DIRECTION INPUT ;
    ANTENNADIFFAREA 1.672500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 4.000 4.500 5.300 ;
        RECT 4.150 3.700 4.650 4.000 ;
        RECT 4.250 1.050 4.500 3.700 ;
      LAYER Metal2 ;
        RECT 4.200 4.000 4.600 4.050 ;
        RECT 4.200 3.700 4.650 4.000 ;
        RECT 4.200 3.650 4.600 3.700 ;
    END
  END X2
  PIN X3
    DIRECTION INPUT ;
    ANTENNADIFFAREA 1.290000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.000 2.600 5.300 ;
        RECT 2.250 1.050 2.500 5.000 ;
      LAYER Metal2 ;
        RECT 2.150 5.300 2.550 5.350 ;
        RECT 2.150 5.000 2.600 5.300 ;
        RECT 2.150 4.950 2.550 5.000 ;
    END
  END X3
  OBS
      LAYER Metal1 ;
        RECT -0.200 2.650 0.050 5.300 ;
        RECT 1.400 3.450 1.650 5.300 ;
        RECT 3.000 5.000 3.500 5.300 ;
        RECT 1.400 2.950 1.900 3.450 ;
        RECT -0.300 2.550 0.200 2.650 ;
        RECT -0.300 2.250 0.300 2.550 ;
        RECT -0.300 2.150 0.200 2.250 ;
        RECT -0.300 1.050 -0.050 2.150 ;
        RECT 1.400 1.050 1.650 2.950 ;
        RECT 3.100 1.050 3.350 5.000 ;
        RECT 5.950 1.250 6.200 5.300 ;
        RECT 7.800 5.000 8.300 5.300 ;
        RECT 5.850 0.950 6.350 1.250 ;
        RECT 7.950 1.050 8.200 5.000 ;
        RECT 9.800 3.150 10.050 5.300 ;
        RECT 9.800 2.900 10.200 3.150 ;
        RECT 9.400 2.150 9.700 2.650 ;
        RECT 9.950 1.250 10.200 2.900 ;
        RECT 9.800 0.950 10.300 1.250 ;
      LAYER Metal2 ;
        RECT 3.050 5.300 3.450 5.350 ;
        RECT 7.850 5.300 8.250 5.350 ;
        RECT 3.050 5.000 8.300 5.300 ;
        RECT 3.050 4.950 3.450 5.000 ;
        RECT 7.850 4.950 8.250 5.000 ;
        RECT -0.150 2.550 0.250 2.600 ;
        RECT 9.350 2.550 9.750 2.600 ;
        RECT -0.200 2.250 9.800 2.550 ;
        RECT -0.150 2.200 0.250 2.250 ;
        RECT 9.300 2.200 9.800 2.250 ;
        RECT 5.900 1.250 6.300 1.300 ;
        RECT 9.850 1.250 10.250 1.300 ;
        RECT 5.900 0.950 10.300 1.250 ;
        RECT 5.900 0.900 6.300 0.950 ;
        RECT 9.850 0.900 10.250 0.950 ;
  END
END gf180mcu_osu_sc_gp9t3v3__mux4_1
END LIBRARY

