* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__mux4_1 VDD C1 C0 VSS X0 X1 OUT X2 X3
X0 a_1160_210# C1 OUT VDD pfet_03v3 ad=0.85p pd=4.4u as=0.595p ps=2.4u w=1.7u l=0.3u
X1 X2 a_250_210# a_590_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 X0 a_250_210# a_1160_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.32p ps=1.65u w=0.85u l=0.3u
X3 X2 C0 a_590_210# VDD pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X4 a_n90_210# C1 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 X0 C0 a_1160_210# VDD pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X6 a_250_210# C0 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 OUT C1 a_590_210# VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 a_n90_210# C1 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_250_210# C0 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X10 OUT a_n90_210# a_590_210# VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X11 a_590_210# C0 X3 VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# C0 X1 VSS nfet_03v3 ad=0.32p pd=1.65u as=0.425p ps=2.7u w=0.85u l=0.3u
X13 a_590_210# a_250_210# X3 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X14 a_1160_210# a_n90_210# OUT VSS nfet_03v3 ad=0.6025p pd=3.2u as=0.2975p ps=1.55u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# X1 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
C0 a_n90_210# OUT 0.1469f
C1 a_250_210# a_590_210# 0.03014f
C2 a_250_210# a_n90_210# 0.08868f
C3 C1 C0 0.05224f
C4 C0 X0 0.08405f
C5 C1 a_1160_210# 0.53587f
C6 X1 a_590_210# 0.03496f
C7 C0 OUT 0.00857f
C8 a_1160_210# X0 0.20363f
C9 C1 VDD 0.4296f
C10 X0 VDD 0.06464f
C11 a_1160_210# OUT 0.22347f
C12 X1 a_n90_210# 0.01914f
C13 a_250_210# C0 0.3665f
C14 OUT VDD 0.05981f
C15 C1 X3 0.01769f
C16 a_250_210# a_1160_210# 0.02157f
C17 X2 C1 0.01928f
C18 a_250_210# VDD 0.90082f
C19 X3 OUT 0
C20 X2 OUT 0
C21 a_250_210# X3 0.37991f
C22 C0 X1 0.06472f
C23 X2 a_250_210# 0.03943f
C24 a_1160_210# X1 0.32933f
C25 X1 VDD 0.05717f
C26 X2 X1 0.37197f
C27 a_n90_210# a_590_210# 0.10428f
C28 C1 X0 0.02056f
C29 C0 a_590_210# 0.25009f
C30 C1 OUT 0.07582f
C31 a_1160_210# a_590_210# 0.03595f
C32 X0 OUT 0.00299f
C33 C0 a_n90_210# 0.52899f
C34 a_590_210# VDD 0.28422f
C35 a_250_210# C1 0.02971f
C36 a_1160_210# a_n90_210# 0.14845f
C37 a_250_210# X0 0.00583f
C38 a_n90_210# VDD 0.51226f
C39 a_250_210# OUT 0
C40 X3 a_590_210# 0.35452f
C41 X2 a_590_210# 0.22961f
C42 X3 a_n90_210# 0.01961f
C43 X2 a_n90_210# 0.02067f
C44 C1 X1 0.01724f
C45 X1 X0 0.01083f
C46 C0 a_1160_210# 0.16894f
C47 C0 VDD 0.41628f
C48 X1 OUT 0
C49 a_1160_210# VDD 0.11048f
C50 a_250_210# X1 0.04064f
C51 C0 X3 0.04882f
C52 X2 C0 0.1344f
C53 a_1160_210# X3 0
C54 X2 a_1160_210# 0.00111f
C55 X3 VDD 0.09082f
C56 X2 VDD 0.06601f
C57 X2 X3 0.0012f
C58 C1 a_590_210# 0.04739f
C59 X0 a_590_210# 0.37242f
C60 a_590_210# OUT 0.34464f
C61 C1 a_n90_210# 1.09377f
C62 a_n90_210# X0 0.05962f
C63 OUT VSS 0.12063f
C64 X0 VSS 0.11727f
C65 X1 VSS 0.09987f
C66 X2 VSS 0.11206f
C67 X3 VSS 0.12356f
C68 C0 VSS 1.0511f
C69 C1 VSS 1.3511f
C70 VDD VSS 5.40678f
C71 a_1160_210# VSS 0.72049f
C72 a_590_210# VSS 0.35695f
C73 a_n90_210# VSS 1.23402f
C74 a_250_210# VSS 1.33984f
.ends

