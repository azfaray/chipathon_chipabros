* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.2.ext - technology: gf180mcuC

X0 a_1160_210# C1.t0 OUT.t1 VDD.t3 pfet_03v3 ad=0.85p pd=4.4u as=0.595p ps=2.4u w=1.7u l=0.3u
X1 X2.t1 a_250_210# a_590_210# VSS.t8 nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 X0.t0 a_250_210# a_1160_210# VSS.t7 nfet_03v3 ad=0.5525p pd=3u as=0.32p ps=1.65u w=0.85u l=0.3u
X3 X2.t0 C0.t0 a_590_210# VDD.t0 pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X4 a_n90_210# C1.t1 VSS.t5 VSS.t4 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 X0.t1 C0.t1 a_1160_210# VDD.t7 pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X6 a_250_210# C0.t2 VSS.t1 VSS.t0 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 OUT.t0 C1.t2 a_590_210# VSS.t3 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 a_n90_210# C1.t3 VDD.t2 VDD.t1 pfet_03v3 ad=1.02p pd=4.6u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_250_210# C0.t3 VDD.t9 VDD.t8 pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X10 OUT.t2 a_n90_210# a_590_210# VDD.t4 pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X11 a_590_210# C0.t4 X3.t0 VSS.t9 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# C0.t5 X1.t0 VSS.t2 nfet_03v3 ad=0.32p pd=1.65u as=0.425p ps=2.7u w=0.85u l=0.3u
X13 a_590_210# a_250_210# X3.t1 VDD.t6 pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X14 a_1160_210# a_n90_210# OUT.t3 VSS.t6 nfet_03v3 ad=0.6025p pd=3.2u as=0.2975p ps=1.55u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# X1.t1 VDD.t5 pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
C0 a_1160_210# X3 0
C1 C1 a_1160_210# 0.53587f
C2 OUT C0 0.00857f
C3 X1 a_250_210# 0.04064f
C4 VDD a_250_210# 0.90091f
C5 a_590_210# X2 0.22961f
C6 a_590_210# X3 0.35452f
C7 a_590_210# C1 0.04739f
C8 X0 C0 0.08405f
C9 OUT a_1160_210# 0.22347f
C10 X2 X3 0.0012f
C11 a_n90_210# C0 0.52899f
C12 X2 C1 0.01928f
C13 C1 X3 0.01769f
C14 X1 VDD 0.05717f
C15 X0 a_1160_210# 0.20363f
C16 a_n90_210# a_1160_210# 0.14865f
C17 a_250_210# C0 0.3665f
C18 a_590_210# OUT 0.34464f
C19 X2 OUT 0
C20 OUT X3 0
C21 OUT C1 0.07582f
C22 a_590_210# X0 0.37242f
C23 a_1160_210# a_250_210# 0.02157f
C24 a_590_210# a_n90_210# 0.1043f
C25 X1 C0 0.06472f
C26 VDD C0 0.41628f
C27 X0 C1 0.02056f
C28 X2 a_n90_210# 0.02067f
C29 a_n90_210# X3 0.01961f
C30 a_n90_210# C1 1.09445f
C31 a_590_210# a_250_210# 0.03014f
C32 X1 a_1160_210# 0.32933f
C33 VDD a_1160_210# 0.11137f
C34 X2 a_250_210# 0.03943f
C35 X3 a_250_210# 0.37991f
C36 C1 a_250_210# 0.02971f
C37 X0 OUT 0.00299f
C38 a_n90_210# OUT 0.1469f
C39 X1 a_590_210# 0.03496f
C40 a_590_210# VDD 0.28462f
C41 X1 X2 0.37197f
C42 X2 VDD 0.06601f
C43 X0 a_n90_210# 0.05962f
C44 X1 C1 0.01724f
C45 VDD X3 0.09082f
C46 OUT a_250_210# 0
C47 a_1160_210# C0 0.16894f
C48 VDD C1 0.4429f
C49 X0 a_250_210# 0.00583f
C50 a_n90_210# a_250_210# 0.08779f
C51 a_590_210# C0 0.25009f
C52 X1 OUT 0
C53 OUT VDD 0.05981f
C54 X2 C0 0.1344f
C55 X3 C0 0.04882f
C56 C1 C0 0.05224f
C57 a_590_210# a_1160_210# 0.03595f
C58 X1 X0 0.01083f
C59 X0 VDD 0.06483f
C60 X1 a_n90_210# 0.01914f
C61 a_n90_210# VDD 0.51227f
C62 X2 a_1160_210# 0.00111f
R0 C1.n0 C1.t2 90.406
R1 C1 C1.n0 50.1755
R2 C1.n1 C1.t1 36.5005
R3 C1.n0 C1.t0 34.6755
R4 C1.n1 C1.t3 29.8088
R5 C1 C1.n1 12.5005
R6 OUT.n2 OUT.n1 6.8405
R7 OUT.n3 OUT.n2 4.5005
R8 OUT.n1 OUT.t3 3.1505
R9 OUT.n2 OUT.n0 2.21083
R10 OUT.n1 OUT.t0 2.03874
R11 OUT.n0 OUT.t1 1.7505
R12 OUT.n0 OUT.t2 1.13285
R13 OUT OUT.n3 0.03425
R14 OUT.n3 OUT 0.03425
R15 VDD.t5 VDD.t0 578.125
R16 VDD.t7 VDD.n2 570.312
R17 VDD.t1 VDD.n7 398.438
R18 VDD.t4 VDD.t3 312.5
R19 VDD.t0 VDD.t6 312.5
R20 VDD.n3 VDD.t5 304.688
R21 VDD.n6 VDD.t6 273.438
R22 VDD.t8 VDD.n6 257.812
R23 VDD.t3 VDD.n1 176.863
R24 VDD.n7 VDD.t8 132.812
R25 VDD VDD.t1 98.538
R26 VDD.n2 VDD.n1 12.6005
R27 VDD.n4 VDD.n3 12.6005
R28 VDD.n6 VDD.n5 12.6005
R29 VDD.n7 VDD.n0 12.6005
R30 VDD.n2 VDD.t4 7.813
R31 VDD.n3 VDD.t7 7.813
R32 VDD VDD.t2 3.3014
R33 VDD.n0 VDD.t9 3.29819
R34 VDD.n5 VDD.n4 0.604786
R35 VDD.n4 VDD.n1 0.238357
R36 VDD VDD.n0 0.199786
R37 VDD.n5 VDD.n0 0.161214
R38 X2.n0 X2.t1 10.2785
R39 X2 X2.n0 4.53425
R40 X2.n0 X2.t0 3.72683
R41 VSS.t8 VSS.t2 1908.73
R42 VSS.n2 VSS.t3 1367.06
R43 VSS.n7 VSS.t9 1109.13
R44 VSS.t4 VSS.n8 1057.54
R45 VSS.t3 VSS.t6 1031.75
R46 VSS.t2 VSS.t7 1031.75
R47 VSS.n3 VSS.t8 748.016
R48 VSS.n8 VSS.t0 696.429
R49 VSS.t0 VSS.n7 644.841
R50 VSS.t6 VSS.n1 604.028
R51 VSS.t7 VSS.n2 541.668
R52 VSS VSS.t4 448.892
R53 VSS.n3 VSS.t9 283.731
R54 VSS.n2 VSS.n1 10.4005
R55 VSS.n4 VSS.n3 10.4005
R56 VSS.n7 VSS.n6 10.4005
R57 VSS.n8 VSS.n0 10.4005
R58 VSS.n5 VSS.t1 8.61774
R59 VSS VSS.t5 8.61774
R60 VSS.n4 VSS.n1 0.527643
R61 VSS VSS.n0 0.186929
R62 VSS.n6 VSS.n4 0.174071
R63 VSS.n6 VSS.n5 0.1355
R64 VSS.n5 VSS.n0 0.0326429
R65 X0.n0 X0.t0 10.2785
R66 X0.n1 X0.n0 4.5005
R67 X0.n0 X0.t1 3.72683
R68 X0 X0.n1 0.03425
R69 X0.n1 X0 0.03425
R70 C0.n1 C0.t4 45.6255
R71 C0.n0 C0.t5 45.6255
R72 C0.n3 C0.t2 36.777
R73 C0.n1 C0.t0 30.4172
R74 C0.n0 C0.t1 30.4172
R75 C0.n3 C0.t3 30.0854
R76 C0.n2 C0.n0 13.3212
R77 C0.n4 C0.n3 12.5005
R78 C0.n2 C0.n1 12.5005
R79 C0.n4 C0.n2 0.808357
R80 C0 C0.n4 0.03425
R81 X3.n0 X3.t0 9.37374
R82 X3 X3.n0 4.79525
R83 X3.n0 X3.t1 2.86619
R84 X1.n0 X1.t0 9.16673
R85 X1 X1.n0 4.53425
R86 X1.n0 X1.t1 3.10919
C63 OUT VSS 0.12063f
C64 X0 VSS 0.11707f
C65 X1 VSS 0.09987f
C66 X2 VSS 0.11206f
C67 X3 VSS 0.12356f
C68 C0 VSS 1.0511f
C69 C1 VSS 1.33736f
C70 VDD VSS 5.51811f
C71 a_1160_210# VSS 0.71945f **FLOATING
C72 a_590_210# VSS 0.35653f **FLOATING
C73 a_n90_210# VSS 1.23339f **FLOATING
C74 a_250_210# VSS 1.3408f **FLOATING
