* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__aoi33_1.2.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__aoi33_1 VDD C B A F E D OUT VSS
X0 a_1310_210# F.t0 VSS.t7 VSS.t6 nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 OUT.t2 D.t0 a_1480_210# VSS.t1 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X2 a_1480_210# E.t0 a_1310_210# VSS.t0 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 a_1310_720# F.t1 OUT.t4 VDD.t8 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 a_1310_720# D.t1 OUT.t1 VDD.t1 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 a_1820_210# A.t0 OUT.t3 VSS.t2 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X6 OUT.t0 E.t1 a_1310_720# VDD.t0 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X7 VSS.t5 C.t0 a_1990_210# VSS.t4 nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X8 a_1990_210# B.t0 a_1820_210# VSS.t3 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X9 VDD.t5 A.t1 a_1310_720# VDD.t4 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X10 VDD.t3 C.t1 a_1310_720# VDD.t2 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X11 a_1310_720# B.t1 VDD.t7 VDD.t6 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
C0 E OUT 0.05861f
C1 D a_1480_210# 0.00297f
C2 D a_1310_720# 0.0172f
C3 A a_1310_720# 0.01969f
C4 A B 0.13834f
C5 OUT a_1820_210# 0.00354f
C6 D F 0
C7 A F 0
C8 E a_1310_720# 0.01759f
C9 E F 0.07113f
C10 C OUT 0.10022f
C11 D VDD 0.08675f
C12 A VDD 0.09996f
C13 OUT a_1480_210# 0.00316f
C14 E VDD 0.08723f
C15 E a_1310_210# 0.00297f
C16 OUT a_1310_720# 0.62324f
C17 B OUT 0.09467f
C18 OUT F 0.11804f
C19 C a_1310_720# 0.00167f
C20 OUT a_1990_210# 0.00297f
C21 B C 0.13834f
C22 C F 0
C23 A D 0.06819f
C24 OUT VDD 0.16687f
C25 OUT a_1310_210# 0.00232f
C26 B a_1310_720# 0.02283f
C27 D E 0.13834f
C28 a_1310_720# F 0.00167f
C29 B F 0
C30 C VDD 0.11096f
C31 B a_1990_210# 0.00297f
C32 a_1310_720# VDD 0.72085f
C33 A a_1820_210# 0.00297f
C34 B VDD 0.09805f
C35 D OUT 0.18649f
C36 A OUT 0.1684f
C37 F VDD 0.13074f
R0 F.n0 F.t0 35.7401
R1 F.n0 F.t1 29.0484
R2 F F.n0 12.5342
R3 VSS.t3 VSS.t2 876.985
R4 VSS.t6 VSS.t0 876.985
R5 VSS.n3 VSS.t4 748.016
R6 VSS.t1 VSS.n6 644.841
R7 VSS.n7 VSS.t1 593.255
R8 VSS.t4 VSS.n2 500.486
R9 VSS.t0 VSS.n7 283.731
R10 VSS.n6 VSS.t2 232.143
R11 VSS.n3 VSS.t3 128.969
R12 VSS.n8 VSS.t6 82.5815
R13 VSS.n4 VSS.n3 10.4005
R14 VSS.n6 VSS.n5 10.4005
R15 VSS.n7 VSS.n0 10.4005
R16 VSS VSS.t7 8.64666
R17 VSS.n2 VSS.t5 8.61774
R18 VSS.n9 VSS.n8 5.2005
R19 VSS.n8 VSS.n1 1.94494
R20 VSS.n5 VSS.n4 0.154786
R21 VSS.n5 VSS.n0 0.154786
R22 VSS.n9 VSS.n0 0.154786
R23 VSS.n4 VSS.n2 0.148357
R24 VSS VSS.n9 0.0165714
R25 D.n0 D.t1 45.6255
R26 D.n0 D.t0 20.6838
R27 D D.n0 12.5342
R28 OUT.n3 OUT.n0 6.8315
R29 OUT.n5 OUT.n4 4.5455
R30 OUT.n2 OUT.t4 3.57419
R31 OUT.n2 OUT.n1 2.7085
R32 OUT.n0 OUT.t3 2.03874
R33 OUT.n0 OUT.t2 2.03874
R34 OUT.n1 OUT.t1 1.13285
R35 OUT.n1 OUT.t0 1.13285
R36 OUT.n4 OUT.n3 1.0115
R37 OUT.n3 OUT.n2 0.4505
R38 OUT OUT.n5 0.03425
R39 OUT.n5 OUT 0.03425
R40 E.n0 E.t1 45.6255
R41 E.n0 E.t0 20.6838
R42 E E.n0 12.5342
R43 VDD.t6 VDD.t4 265.625
R44 VDD.t8 VDD.t0 265.625
R45 VDD.n4 VDD.t2 226.562
R46 VDD.t1 VDD.n8 195.312
R47 VDD.n9 VDD.t1 179.689
R48 VDD.t2 VDD.n3 161.044
R49 VDD.t0 VDD.n9 85.938
R50 VDD.n8 VDD.t4 70.313
R51 VDD.n4 VDD.t6 39.063
R52 VDD.n10 VDD.t8 29.738
R53 VDD.n5 VDD.n4 12.6005
R54 VDD.n8 VDD.n7 12.6005
R55 VDD.n9 VDD.n0 12.6005
R56 VDD VDD.n10 6.3005
R57 VDD.n3 VDD.t3 3.29819
R58 VDD.n6 VDD.n2 2.9425
R59 VDD.n10 VDD.n1 1.7505
R60 VDD.n2 VDD.t7 1.13285
R61 VDD.n2 VDD.t5 1.13285
R62 VDD.n7 VDD.n0 0.154786
R63 VDD VDD.n0 0.154786
R64 VDD.n5 VDD.n3 0.148357
R65 VDD.n7 VDD.n6 0.0840714
R66 VDD.n6 VDD.n5 0.0712143
R67 A.n0 A.t1 45.6255
R68 A.n0 A.t0 20.6838
R69 A A.n0 12.5342
R70 C.n0 C.t1 45.6255
R71 C.n0 C.t0 20.6838
R72 C C.n0 12.5342
R73 B.n0 B.t1 45.6255
R74 B.n0 B.t0 20.6838
R75 B B.n0 12.5342
C38 OUT VSS 0.42067f
C39 C VSS 0.39621f
C40 B VSS 0.30452f
C41 A VSS 0.30946f
C42 D VSS 0.30954f
C43 E VSS 0.32807f
C44 F VSS 0.39864f
C45 VDD VSS 2.97769f
C46 a_1990_210# VSS 0.00795f **FLOATING
C47 a_1820_210# VSS 0.00738f **FLOATING
C48 a_1480_210# VSS 0.00738f **FLOATING
C49 a_1310_210# VSS 0.00795f **FLOATING
C50 a_1310_720# VSS 0.07075f **FLOATING
.ends gf180mcu_osu_sc_gp9t3v3__aoi33_1
