* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.ext - technology: gf180mcuD

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

.subckt gf180mcu_osu_sc_gp9t3v3__mux4_1 VDD C1 C0 VSS X0 X1 OUT X2 X3
X0 a_1160_210# C1 OUT VDD pfet_03v3 ad=0.85p pd=4.4u as=0.595p ps=2.4u w=1.7u l=0.3u
X1 X2 a_250_210# a_590_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 X0 a_250_210# a_1160_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.32p ps=1.65u w=0.85u l=0.3u
X3 X2 C0 a_590_210# VDD pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X4 a_n90_210# C1 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 X0 C0 a_1160_210# VDD pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X6 a_250_210# C0 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 OUT C1 a_590_210# VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 a_n90_210# C1 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_250_210# C0 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X10 OUT a_n90_210# a_590_210# VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X11 a_590_210# C0 X3 VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# C0 X1 VSS nfet_03v3 ad=0.32p pd=1.65u as=0.425p ps=2.7u w=0.85u l=0.3u
X13 a_590_210# a_250_210# X3 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X14 a_1160_210# a_n90_210# OUT VSS nfet_03v3 ad=0.6025p pd=3.2u as=0.2975p ps=1.55u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# X1 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
.ends gf180mcu_osu_sc_gp9t3v3__mux4_1


VDD VDD 0 3.3
VSS VSS 0 0

VC0 C0 0 PULSE(0 3.3 0ns 0.5ns 0.5ns 19.98ns 40ns)
VC1 C1 0 PULSE(0 3.3 0ns 0.5ns 0.5ns 39.98ns 80ns)

VX0 X0 0 PULSE(0 3.3 0ns 0.5ns 0.5ns 9.98ns 20ns)
VX1 X1 0 PULSE(0 3.3 0ns 0.5ns 0.5ns 4.98ns 10ns)
VX2 X2 0 3.3
VX3 X3 0 0

* DUT
Xdut VDD C1 C0 VSS X0 X1 OUT X2 X3 gf180mcu_osu_sc_gp9t3v3__mux4_1


* Simulation
.tran 0.1n 100n

.control

run
set color0=white
set color1=black
set xbrushwidth=3
plot out x0+4 x1+8 x2+12 x3+16 C0+20 C1+24
.endc

.end
