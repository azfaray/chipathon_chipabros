* tb_aoi33.spice  — AOI33 extracted cell functional check

* --- GF180MCU-D models (your lines) ---
.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib     /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

.subckt gf180mcu_osu_sc_gp9t3v3__aoi33_1 F E D A B C OUT VDD VSS
X0 a_1310_210# F VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 OUT D a_1480_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X2 a_1480_210# E a_1310_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 a_1310_720# F OUT VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 a_1310_720# D OUT VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 a_1820_210# A OUT VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X6 OUT E a_1310_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X7 VSS C a_1990_210# VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X8 a_1990_210# B a_1820_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X9 VDD A a_1310_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X10 VDD C a_1310_720# VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X11 a_1310_720# B VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
.ends

VDD VDD 0 3.3
VSS VSS 0 0

.param T0=50n tr=2n tf=2n
VA A 0  PULSE(0 3.3 0 {tr} {tf} {T0/2}   {T0})
VB B 0  PULSE(0 3.3 0 {tr} {tf} {T0}     {2*T0})
VC C 0  PULSE(0 3.3 0 {tr} {tf} {2*T0}   {4*T0})
VD D 0  PULSE(0 3.3 0 {tr} {tf} {4*T0}   {8*T0})
VE E 0  PULSE(0 3.3 0 {tr} {tf} {8*T0}   {16*T0})
VF F 0  PULSE(0 3.3 0 {tr} {tf} {16*T0}  {32*T0})

* --- DUT + load (mind the pin order: F E D A B C OUT VDD VSS) ---
XU1 F E D A B C OUT VDD VSS gf180mcu_osu_sc_gp9t3v3__aoi33_1
Cload OUT 0 10f


.tran 50n {32*T0}
.control
  set color0=white
  set color1=black
  set linewidth=5
  run
  setplot tran1
  plot v(out) v(a)+4 v(b)+8 v(c)+12 v(d)+16 v(e)+20 v(f)+24
.endc
.end
