* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.2.ext - technology: gf180mcuC

X0 a_1160_210# C1.t0 OUT.t3 VDD.t3 pfet_03v3 ad=0.85p pd=4.4u as=0.595p ps=2.4u w=1.7u l=0.3u
X1 X2.t0 a_250_210# a_590_210# VSS.t7 nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 X0.t1 a_250_210# a_1160_210# VSS.t6 nfet_03v3 ad=0.5525p pd=3u as=0.32p ps=1.65u w=0.85u l=0.3u
X3 X2.t1 C0.t0 a_590_210# VDD.t9 pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X4 a_n90_210# C1.t1 VSS.t3 VSS.t2 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 X0.t0 C0.t1 a_1160_210# VDD.t4 pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X6 a_250_210# C0.t2 VSS.t5 VSS.t4 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 OUT.t2 C1.t2 a_590_210# VSS.t1 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 a_n90_210# C1.t3 VDD.t2 VDD.t1 pfet_03v3 ad=1.02p pd=4.6u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_250_210# C0.t3 VDD.t6 VDD.t5 pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X10 OUT.t0 a_n90_210# a_590_210# VDD.t0 pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X11 a_590_210# C0.t4 X3.t0 VSS.t9 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# C0.t5 X1.t0 VSS.t8 nfet_03v3 ad=0.32p pd=1.65u as=0.425p ps=2.7u w=0.85u l=0.3u
X13 a_590_210# a_250_210# X3.t1 VDD.t8 pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X14 a_1160_210# a_n90_210# OUT.t1 VSS.t0 nfet_03v3 ad=0.6025p pd=3.2u as=0.2975p ps=1.55u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# X1.t1 VDD.t7 pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
C0 OUT C0 0.00857f
C1 a_250_210# a_n90_210# 0.08868f
C2 a_590_210# X2 0.22961f
C3 C0 a_n90_210# 0.52899f
C4 X3 VDD 0.09082f
C5 C1 VDD 0.4296f
C6 a_590_210# X1 0.03496f
C7 X0 X1 0.01083f
C8 OUT X3 0
C9 X2 VDD 0.06601f
C10 OUT C1 0.07582f
C11 a_250_210# a_1160_210# 0.02157f
C12 X3 a_n90_210# 0.01961f
C13 a_1160_210# C0 0.16894f
C14 a_n90_210# C1 1.09377f
C15 OUT X2 0
C16 X1 VDD 0.05717f
C17 a_n90_210# X2 0.02067f
C18 a_590_210# X0 0.37242f
C19 a_250_210# C0 0.3665f
C20 OUT X1 0
C21 X3 a_1160_210# 0
C22 a_n90_210# X1 0.01914f
C23 a_1160_210# C1 0.53587f
C24 a_590_210# VDD 0.28422f
C25 X0 VDD 0.06464f
C26 a_1160_210# X2 0.00111f
C27 X3 a_250_210# 0.37991f
C28 OUT a_590_210# 0.34464f
C29 OUT X0 0.00299f
C30 X3 C0 0.04882f
C31 a_250_210# C1 0.02971f
C32 C0 C1 0.05224f
C33 a_590_210# a_n90_210# 0.10428f
C34 a_n90_210# X0 0.05962f
C35 a_1160_210# X1 0.32933f
C36 a_250_210# X2 0.03943f
C37 C0 X2 0.1344f
C38 OUT VDD 0.05981f
C39 a_250_210# X1 0.04064f
C40 a_n90_210# VDD 0.51226f
C41 X3 C1 0.01769f
C42 C0 X1 0.06472f
C43 a_1160_210# a_590_210# 0.03595f
C44 a_1160_210# X0 0.20363f
C45 X3 X2 0.0012f
C46 OUT a_n90_210# 0.1469f
C47 X2 C1 0.01928f
C48 a_250_210# a_590_210# 0.03014f
C49 a_250_210# X0 0.00583f
C50 a_1160_210# VDD 0.11048f
C51 a_590_210# C0 0.25009f
C52 C0 X0 0.08405f
C53 X1 C1 0.01724f
C54 OUT a_1160_210# 0.22347f
C55 X2 X1 0.37197f
C56 a_250_210# VDD 0.90082f
C57 a_1160_210# a_n90_210# 0.14845f
C58 C0 VDD 0.41628f
C59 X3 a_590_210# 0.35452f
C60 OUT a_250_210# 0
C61 a_590_210# C1 0.04739f
C62 X0 C1 0.02056f
R0 C1.n0 C1.t2 90.406
R1 C1 C1.n0 50.1755
R2 C1.n1 C1.t1 36.5005
R3 C1.n0 C1.t0 34.6755
R4 C1.n1 C1.t3 29.8088
R5 C1 C1.n1 12.5005
R6 OUT.n2 OUT.n1 6.8405
R7 OUT.n3 OUT.n2 4.5005
R8 OUT.n1 OUT.t1 3.1505
R9 OUT.n2 OUT.n0 2.21083
R10 OUT.n1 OUT.t2 2.03874
R11 OUT.n0 OUT.t3 1.7505
R12 OUT.n0 OUT.t0 1.13285
R13 OUT OUT.n3 0.03425
R14 OUT.n3 OUT 0.03425
R15 VDD.t7 VDD.t9 578.125
R16 VDD.t4 VDD.n2 570.312
R17 VDD.t1 VDD.n7 398.438
R18 VDD.t0 VDD.t3 312.5
R19 VDD.t9 VDD.t8 312.5
R20 VDD.n3 VDD.t7 304.688
R21 VDD.n6 VDD.t8 273.438
R22 VDD.t5 VDD.n6 257.812
R23 VDD.t3 VDD.n1 176.863
R24 VDD.n7 VDD.t5 132.812
R25 VDD VDD.t1 98.538
R26 VDD.n2 VDD.n1 12.6005
R27 VDD.n4 VDD.n3 12.6005
R28 VDD.n6 VDD.n5 12.6005
R29 VDD.n7 VDD.n0 12.6005
R30 VDD.n2 VDD.t0 7.813
R31 VDD.n3 VDD.t4 7.813
R32 VDD VDD.t2 3.3014
R33 VDD.n0 VDD.t6 3.29819
R34 VDD.n5 VDD.n4 0.604786
R35 VDD.n4 VDD.n1 0.238357
R36 VDD VDD.n0 0.199786
R37 VDD.n5 VDD.n0 0.161214
R38 X2.n0 X2.t0 10.2785
R39 X2 X2.n0 4.53425
R40 X2.n0 X2.t1 3.72683
R41 VSS.t7 VSS.t8 1908.73
R42 VSS.n2 VSS.t1 1367.06
R43 VSS.t2 VSS.n7 1315.48
R44 VSS.t1 VSS.t0 1031.75
R45 VSS.t8 VSS.t6 1031.75
R46 VSS.t4 VSS.n6 902.779
R47 VSS.n6 VSS.t9 851.191
R48 VSS.n3 VSS.t7 748.016
R49 VSS.t0 VSS.n1 604.028
R50 VSS.t6 VSS.n2 541.668
R51 VSS VSS.t2 448.892
R52 VSS.n7 VSS.t4 438.493
R53 VSS.n3 VSS.t9 283.731
R54 VSS.n2 VSS.n1 10.4005
R55 VSS.n4 VSS.n3 10.4005
R56 VSS.n6 VSS.n5 10.4005
R57 VSS.n7 VSS.n0 10.4005
R58 VSS.n0 VSS.t5 8.61774
R59 VSS VSS.t3 8.61774
R60 VSS.n4 VSS.n1 0.527643
R61 VSS VSS.n0 0.219071
R62 VSS.n5 VSS.n0 0.167643
R63 VSS.n5 VSS.n4 0.141929
R64 X0.n0 X0.t1 10.2785
R65 X0.n1 X0.n0 4.5005
R66 X0.n0 X0.t0 3.72683
R67 X0 X0.n1 0.03425
R68 X0.n1 X0 0.03425
R69 C0.n1 C0.t4 45.6255
R70 C0.n0 C0.t5 45.6255
R71 C0.n3 C0.t2 36.777
R72 C0.n1 C0.t0 30.4172
R73 C0.n0 C0.t1 30.4172
R74 C0.n3 C0.t3 30.0854
R75 C0.n2 C0.n0 13.3212
R76 C0.n4 C0.n3 12.5005
R77 C0.n2 C0.n1 12.5005
R78 C0.n4 C0.n2 0.808357
R79 C0 C0.n4 0.03425
R80 X3.n0 X3.t0 9.37374
R81 X3 X3.n0 4.79525
R82 X3.n0 X3.t1 2.86619
R83 X1.n0 X1.t0 9.16673
R84 X1 X1.n0 4.53425
R85 X1.n0 X1.t1 3.10919
C63 OUT VSS 0.12063f
C64 X0 VSS 0.11727f
C65 X1 VSS 0.09987f
C66 X2 VSS 0.11206f
C67 X3 VSS 0.12356f
C68 C0 VSS 1.0511f
C69 C1 VSS 1.3511f
C70 VDD VSS 5.40678f
C71 a_1160_210# VSS 0.72049f **FLOATING
C72 a_590_210# VSS 0.35695f **FLOATING
C73 a_n90_210# VSS 1.23402f **FLOATING
C74 a_250_210# VSS 1.33984f **FLOATING
