magic
tech gf180mcuC
timestamp 1756902939
<< nwell >>
rect -34 63 215 127
<< nmos >>
rect -15 21 -9 38
rect 19 21 25 38
rect 53 21 59 38
rect 73 21 79 38
rect 110 21 116 38
rect 130 21 136 38
rect 167 21 173 38
rect 187 21 193 38
<< pmos >>
rect -15 72 -9 106
rect 19 72 25 106
rect 53 72 59 106
rect 73 72 79 106
rect 110 72 116 106
rect 130 72 136 106
rect 167 72 173 106
rect 187 72 193 106
<< ndiff >>
rect -25 36 -15 38
rect -25 23 -23 36
rect -18 23 -15 36
rect -25 21 -15 23
rect -9 36 1 38
rect -9 23 -6 36
rect -1 23 1 36
rect -9 21 1 23
rect 9 36 19 38
rect 9 23 11 36
rect 16 23 19 36
rect 9 21 19 23
rect 25 36 35 38
rect 25 23 28 36
rect 33 23 35 36
rect 25 21 35 23
rect 43 36 53 38
rect 43 23 45 36
rect 50 23 53 36
rect 43 21 53 23
rect 59 36 73 38
rect 59 23 62 36
rect 67 23 73 36
rect 59 21 73 23
rect 79 36 92 38
rect 79 23 85 36
rect 90 23 92 36
rect 79 21 92 23
rect 100 36 110 38
rect 100 23 102 36
rect 107 23 110 36
rect 100 21 110 23
rect 116 36 130 38
rect 116 25 119 36
rect 124 25 130 36
rect 116 21 130 25
rect 136 36 149 38
rect 136 23 142 36
rect 147 23 149 36
rect 136 21 149 23
rect 118 19 127 21
rect 157 36 167 38
rect 157 23 159 36
rect 164 23 167 36
rect 157 21 167 23
rect 173 36 187 38
rect 173 23 176 36
rect 181 23 187 36
rect 173 21 187 23
rect 193 36 206 38
rect 193 25 199 36
rect 204 25 206 36
rect 193 21 206 25
rect 196 19 206 21
<< pdiff >>
rect -25 104 -15 106
rect -25 74 -23 104
rect -18 74 -15 104
rect -25 72 -15 74
rect -9 104 3 106
rect -9 74 -4 104
rect 1 74 3 104
rect -9 72 3 74
rect 9 104 19 106
rect 9 74 11 104
rect 16 74 19 104
rect 9 72 19 74
rect 25 104 35 106
rect 25 74 28 104
rect 33 74 35 104
rect 42 100 53 106
rect 25 72 35 74
rect 43 74 45 100
rect 50 74 53 100
rect 43 72 53 74
rect 59 100 73 106
rect 59 74 62 100
rect 67 74 73 100
rect 59 72 73 74
rect 79 104 92 106
rect 79 80 85 104
rect 90 80 92 104
rect 100 104 110 106
rect 100 80 102 104
rect 107 80 110 104
rect 79 74 93 80
rect 99 74 110 80
rect 79 72 92 74
rect 100 72 110 74
rect 116 104 130 106
rect 116 74 119 104
rect 124 74 130 104
rect 116 72 130 74
rect 136 104 149 106
rect 136 80 142 104
rect 147 80 149 104
rect 156 100 167 106
rect 136 74 150 80
rect 157 74 159 100
rect 164 74 167 100
rect 136 72 149 74
rect 157 72 167 74
rect 173 104 187 106
rect 173 74 176 104
rect 181 74 187 104
rect 173 72 187 74
rect 193 104 203 106
rect 193 74 196 104
rect 201 74 203 104
rect 193 72 203 74
<< ndiffc >>
rect -23 23 -18 36
rect -6 23 -1 36
rect 11 23 16 36
rect 28 23 33 36
rect 45 23 50 36
rect 62 23 67 36
rect 85 23 90 36
rect 102 23 107 36
rect 119 25 124 36
rect 142 23 147 36
rect 159 23 164 36
rect 176 23 181 36
rect 199 25 204 36
<< pdiffc >>
rect -23 74 -18 104
rect -4 74 1 104
rect 11 74 16 104
rect 28 74 33 104
rect 45 74 50 100
rect 62 74 67 100
rect 85 80 90 104
rect 102 80 107 104
rect 119 74 124 104
rect 142 80 147 104
rect 159 74 164 100
rect 176 74 181 104
rect 196 74 201 104
<< psubdiff >>
rect -26 11 -15 13
rect -26 6 -23 11
rect -18 6 -15 11
rect -26 4 -15 6
rect 8 11 19 13
rect 8 6 11 11
rect 16 6 19 11
rect 8 4 19 6
rect 34 11 45 13
rect 34 6 37 11
rect 42 6 45 11
rect 34 4 45 6
rect 56 11 67 13
rect 56 6 59 11
rect 64 6 67 11
rect 138 11 149 13
rect 56 4 67 6
rect 138 6 141 11
rect 146 6 149 11
rect 196 11 207 13
rect 138 4 149 6
rect 196 6 199 11
rect 204 6 207 11
rect 196 4 207 6
<< nsubdiff >>
rect -26 120 -15 122
rect -26 115 -23 120
rect -18 115 -15 120
rect -26 113 -15 115
rect 8 120 19 122
rect 8 115 11 120
rect 16 115 19 120
rect 8 113 19 115
rect 33 120 44 122
rect 127 120 138 122
rect 33 115 36 120
rect 41 115 44 120
rect 33 113 44 115
rect 127 115 130 120
rect 135 115 138 120
rect 127 113 138 115
rect 164 120 175 122
rect 164 115 167 120
rect 172 115 175 120
rect 164 113 175 115
rect 195 120 206 122
rect 195 115 198 120
rect 203 115 206 120
rect 195 113 206 115
<< psubdiffcont >>
rect -23 6 -18 11
rect 11 6 16 11
rect 37 6 42 11
rect 59 6 64 11
rect 141 6 146 11
rect 199 6 204 11
<< nsubdiffcont >>
rect -23 115 -18 120
rect 11 115 16 120
rect 36 115 41 120
rect 130 115 135 120
rect 167 115 172 120
rect 198 115 203 120
<< polysilicon >>
rect 53 116 116 120
rect -15 106 -9 111
rect 19 106 25 111
rect 53 106 59 116
rect 73 106 79 111
rect 110 106 116 116
rect 130 106 136 111
rect 167 106 173 111
rect 187 106 193 111
rect 205 75 215 77
rect -15 67 -9 72
rect 19 67 25 72
rect 53 69 59 72
rect -21 65 -9 67
rect -21 59 -19 65
rect -13 59 -9 65
rect -21 57 -9 59
rect 14 65 25 67
rect 14 59 16 65
rect 22 59 25 65
rect 30 67 59 69
rect 73 67 79 72
rect 110 69 116 72
rect 30 61 32 67
rect 38 64 59 67
rect 70 65 80 67
rect 38 61 40 64
rect 30 59 40 61
rect 70 60 72 65
rect 62 59 72 60
rect 78 59 80 65
rect 14 57 25 59
rect -15 38 -9 57
rect 19 38 25 57
rect 62 56 80 59
rect 94 65 116 69
rect 130 67 136 72
rect 167 70 173 72
rect 127 65 137 67
rect 62 49 68 56
rect 94 51 100 65
rect 127 60 129 65
rect 53 44 68 49
rect 73 46 100 51
rect 119 59 129 60
rect 135 59 137 65
rect 119 56 137 59
rect 151 65 173 70
rect 119 50 125 56
rect 53 38 59 44
rect 73 38 79 46
rect 110 45 125 50
rect 110 38 116 45
rect 130 38 136 45
rect -15 15 -9 21
rect 19 16 25 21
rect 53 16 59 21
rect 73 11 79 21
rect 110 16 116 21
rect 130 11 136 21
rect 73 7 136 11
rect 151 11 155 65
rect 187 63 193 72
rect 205 69 207 75
rect 213 69 215 75
rect 205 67 215 69
rect 183 62 198 63
rect 207 62 213 67
rect 178 61 213 62
rect 176 60 213 61
rect 175 58 213 60
rect 175 57 183 58
rect 199 57 213 58
rect 175 49 181 57
rect 167 44 181 49
rect 186 51 196 53
rect 186 45 188 51
rect 194 45 196 51
rect 167 38 173 44
rect 186 43 196 45
rect 187 38 193 43
rect 167 16 173 21
rect 187 11 193 21
rect 151 7 193 11
<< polycontact >>
rect -19 59 -13 65
rect 16 59 22 65
rect 32 61 38 67
rect 72 59 78 65
rect 129 59 135 65
rect 207 69 213 75
rect 188 45 194 51
<< metal1 >>
rect -34 120 215 127
rect -34 115 -23 120
rect -18 115 11 120
rect 16 115 36 120
rect 41 115 130 120
rect 135 115 167 120
rect 172 115 198 120
rect 203 115 215 120
rect -34 113 215 115
rect -23 104 -18 113
rect -23 72 -18 74
rect -4 104 1 106
rect -21 59 -19 65
rect -13 59 -11 65
rect -4 53 1 74
rect 11 104 16 113
rect 11 72 16 74
rect 28 104 33 106
rect 42 100 44 106
rect 50 100 52 106
rect 60 100 62 106
rect 68 100 70 106
rect 85 104 90 106
rect 28 69 33 74
rect 28 67 38 69
rect 16 65 22 67
rect 16 57 22 59
rect 28 61 32 67
rect 28 59 38 61
rect -6 51 4 53
rect -6 45 -2 51
rect 4 45 6 51
rect -6 43 4 45
rect -23 36 -18 38
rect -23 14 -18 23
rect -6 36 -1 43
rect -6 21 -1 23
rect 11 36 16 38
rect 11 14 16 23
rect 28 36 33 59
rect 28 21 33 23
rect 45 36 50 74
rect 45 21 50 23
rect 102 104 107 106
rect 119 104 124 106
rect 83 74 85 80
rect 91 74 93 80
rect 99 74 101 80
rect 107 74 109 80
rect 142 104 147 106
rect 156 100 158 106
rect 164 100 166 106
rect 176 104 181 106
rect 140 74 142 80
rect 148 74 150 80
rect 62 36 67 74
rect 72 65 78 67
rect 72 57 78 59
rect 62 21 67 23
rect 85 36 90 74
rect 85 21 90 23
rect 102 36 107 74
rect 119 36 124 74
rect 129 65 135 67
rect 129 57 135 59
rect 142 36 147 74
rect 102 21 107 23
rect 117 19 119 25
rect 125 19 127 25
rect 142 21 147 23
rect 159 36 164 74
rect 176 64 181 74
rect 171 58 173 64
rect 179 58 181 64
rect 196 104 201 106
rect 196 63 201 74
rect 207 75 213 77
rect 207 67 213 69
rect 196 58 204 63
rect 159 21 164 23
rect 176 36 181 58
rect 188 51 194 53
rect 188 43 194 45
rect 199 36 204 58
rect 176 21 181 23
rect 196 19 198 25
rect 204 19 206 25
rect -34 11 215 14
rect -34 6 -23 11
rect -18 6 11 11
rect 16 6 37 11
rect 42 6 59 11
rect 64 6 141 11
rect 146 6 199 11
rect 204 6 215 11
rect -34 0 215 6
<< via1 >>
rect -19 59 -13 65
rect 44 100 50 106
rect 62 100 68 106
rect 16 59 22 65
rect -2 45 4 51
rect 85 74 91 80
rect 101 74 107 80
rect 158 100 164 106
rect 142 74 148 80
rect 72 59 78 65
rect 129 59 135 65
rect 119 19 125 25
rect 173 58 179 64
rect 207 69 213 75
rect 188 45 194 51
rect 198 19 204 25
<< metal2 >>
rect 43 106 51 107
rect 61 106 69 107
rect 157 106 165 107
rect 43 100 44 106
rect 50 100 52 106
rect 61 100 62 106
rect 68 100 158 106
rect 164 100 166 106
rect 43 99 51 100
rect 61 99 69 100
rect 157 99 165 100
rect 84 80 92 81
rect 100 80 108 81
rect 141 80 149 81
rect 84 74 85 80
rect 91 74 93 80
rect 100 74 101 80
rect 107 74 109 80
rect 141 74 142 80
rect 148 74 150 80
rect 206 75 214 76
rect 84 73 92 74
rect 100 73 108 74
rect 141 73 149 74
rect 206 69 207 75
rect 213 69 214 75
rect 206 68 214 69
rect -20 65 -12 66
rect 15 65 23 66
rect 70 65 80 66
rect 127 65 137 66
rect -20 59 -19 65
rect -13 59 -11 65
rect 15 59 16 65
rect 22 59 72 65
rect 78 59 129 65
rect 135 59 137 65
rect 172 64 181 65
rect -20 38 -12 59
rect 15 58 23 59
rect 71 58 79 59
rect 128 58 136 59
rect 172 58 173 64
rect 179 58 181 64
rect 172 57 181 58
rect -3 51 5 52
rect 187 51 195 52
rect -4 45 -2 51
rect 4 45 188 51
rect 194 45 196 51
rect -3 44 5 45
rect 186 44 196 45
rect 207 38 213 68
rect -20 32 213 38
rect 118 25 126 26
rect 197 25 205 26
rect 118 19 119 25
rect 125 19 198 25
rect 204 19 206 25
rect 118 18 126 19
rect 197 18 205 19
<< labels >>
rlabel metal1 -23 115 -18 120 1 VDD
port 1 n default bidirectional
rlabel metal2 -19 59 -13 65 7 C1
port 2 w default input
rlabel metal2 16 59 22 65 7 C0
port 3 w default input
rlabel metal1 -23 6 -18 11 5 VSS
port 4 s default bidirectional
rlabel metal2 142 74 148 80 3 X0
port 5 e default input
rlabel metal2 101 74 107 80 0 X1
port 6 nsew default input
rlabel metal2 173 58 179 64 3 OUT
port 7 e default output
rlabel metal2 85 74 91 80 0 X2
port 8 nsew default input
rlabel metal2 44 100 50 106 7 X3
port 9 w default input
<< end >>
