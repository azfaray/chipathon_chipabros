* NGSPICE file created from MUX4.ext - technology: gf180mcuC

.subckt MUX4 OUT X0 X1 X3 X2 C1 C0 VDD VSS
X0 a_1160_210# C1 OUT VDD pfet_03v3 ad=0.85p pd=4.4u as=0.595p ps=2.4u w=1.7u l=0.3u
X1 X2 a_250_210# a_590_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 X0 a_250_210# a_1160_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.32p ps=1.65u w=0.85u l=0.3u
X3 X2 C0 a_590_210# VDD pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X4 a_n90_210# C1 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 X0 C0 a_1160_210# VDD pfet_03v3 ad=1.12p pd=4.8u as=0.595p ps=2.4u w=1.7u l=0.3u
X6 a_250_210# C0 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 OUT C1 a_590_210# VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 a_n90_210# C1 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_250_210# C0 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X10 OUT a_n90_210# a_590_210# VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X11 a_590_210# C0 X3 VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# C0 X1 VSS nfet_03v3 ad=0.32p pd=1.65u as=0.425p ps=2.7u w=0.85u l=0.3u
X13 a_590_210# a_250_210# X3 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
X14 a_1160_210# a_n90_210# OUT VSS nfet_03v3 ad=0.6025p pd=3.2u as=0.2975p ps=1.55u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# X1 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.865p ps=4.5u w=1.7u l=0.3u
.ends

