magic
tech gf180mcuD
timestamp 1755592685
<< nwell >>
rect -16 42 283 95
<< nmos >>
rect 3 -1 9 16
rect 45 -1 51 16
rect 65 -1 71 16
rect 113 -1 119 16
rect 142 -1 148 16
rect 177 -1 183 16
rect 221 -1 227 16
rect 250 -1 256 16
<< pmos >>
rect 3 52 9 86
rect 45 52 51 86
rect 65 52 71 86
rect 113 52 119 86
rect 142 52 148 86
rect 177 52 183 86
rect 221 52 227 86
rect 250 52 256 86
<< ndiff >>
rect -7 9 3 16
rect -7 4 -5 9
rect 0 4 3 9
rect -7 -1 3 4
rect 9 9 19 16
rect 9 4 12 9
rect 17 4 19 9
rect 9 -1 19 4
rect 25 9 45 16
rect 25 4 27 9
rect 32 4 45 9
rect 25 -1 45 4
rect 51 9 65 16
rect 51 4 56 9
rect 61 4 65 9
rect 51 -1 65 4
rect 71 9 84 16
rect 71 4 75 9
rect 80 4 84 9
rect 71 -1 84 4
rect 93 9 113 16
rect 93 4 95 9
rect 100 4 113 9
rect 93 -1 113 4
rect 119 9 142 16
rect 119 4 124 9
rect 129 4 142 9
rect 119 -1 142 4
rect 148 9 161 16
rect 148 2 151 9
rect 158 2 161 9
rect 148 -1 161 2
rect 167 9 177 16
rect 167 4 169 9
rect 174 4 177 9
rect 167 -1 177 4
rect 183 9 193 16
rect 183 4 186 9
rect 191 4 193 9
rect 183 -1 193 4
rect 201 9 221 16
rect 201 4 203 9
rect 208 4 221 9
rect 201 -1 221 4
rect 227 9 250 16
rect 227 4 232 9
rect 237 4 250 9
rect 227 -1 250 4
rect 256 9 269 16
rect 256 4 260 9
rect 265 4 269 9
rect 256 -1 269 4
<< pdiff >>
rect -7 81 3 86
rect -7 76 -5 81
rect 0 76 3 81
rect -7 63 3 76
rect -7 58 -5 63
rect 0 58 3 63
rect -7 52 3 58
rect 9 81 19 86
rect 9 76 12 81
rect 17 76 19 81
rect 9 63 19 76
rect 9 58 12 63
rect 17 58 19 63
rect 9 52 19 58
rect 25 81 45 86
rect 25 76 27 81
rect 36 76 45 81
rect 25 63 45 76
rect 25 58 27 63
rect 32 58 45 63
rect 25 52 45 58
rect 51 81 65 86
rect 51 76 56 81
rect 61 76 65 81
rect 51 63 65 76
rect 51 58 56 63
rect 61 58 65 63
rect 51 52 65 58
rect 71 66 87 86
rect 71 61 77 66
rect 82 61 87 66
rect 71 52 87 61
rect 93 66 113 86
rect 93 61 99 66
rect 104 61 113 66
rect 93 52 113 61
rect 119 67 142 86
rect 119 59 124 67
rect 132 59 142 67
rect 119 52 142 59
rect 148 63 161 86
rect 148 58 152 63
rect 157 58 161 63
rect 148 52 161 58
rect 167 81 177 86
rect 167 76 169 81
rect 174 76 177 81
rect 167 63 177 76
rect 167 58 169 63
rect 174 58 177 63
rect 167 52 177 58
rect 183 81 193 86
rect 183 76 186 81
rect 191 76 193 81
rect 183 63 193 76
rect 183 58 186 63
rect 191 58 193 63
rect 183 52 193 58
rect 201 66 221 86
rect 201 61 207 66
rect 212 61 221 66
rect 201 52 221 61
rect 227 66 250 86
rect 227 61 232 66
rect 240 61 250 66
rect 227 52 250 61
rect 256 82 274 86
rect 256 77 262 82
rect 267 77 274 82
rect 256 52 274 77
<< ndiffc >>
rect -5 4 0 9
rect 12 4 17 9
rect 27 4 32 9
rect 56 4 61 9
rect 75 4 80 9
rect 95 4 100 9
rect 124 4 129 9
rect 151 2 158 9
rect 169 4 174 9
rect 186 4 191 9
rect 203 4 208 9
rect 232 4 237 9
rect 260 4 265 9
<< pdiffc >>
rect -5 76 0 81
rect -5 58 0 63
rect 12 76 17 81
rect 12 58 17 63
rect 27 76 36 81
rect 27 58 32 63
rect 56 76 61 81
rect 56 58 61 63
rect 77 61 82 66
rect 99 61 104 66
rect 124 59 132 67
rect 152 58 157 63
rect 169 76 174 81
rect 169 58 174 63
rect 186 76 191 81
rect 186 58 191 63
rect 207 61 212 66
rect 232 61 240 66
rect 262 77 267 82
<< psubdiff >>
rect -7 -14 2 -12
rect -7 -19 -5 -14
rect 0 -19 2 -14
rect -7 -21 2 -19
rect 12 -14 21 -12
rect 12 -19 14 -14
rect 19 -19 21 -14
rect 12 -21 21 -19
rect 31 -14 40 -12
rect 31 -19 33 -14
rect 38 -19 40 -14
rect 31 -21 40 -19
rect 50 -14 59 -12
rect 50 -19 52 -14
rect 57 -19 59 -14
rect 50 -21 59 -19
rect 69 -14 78 -12
rect 69 -19 71 -14
rect 76 -19 78 -14
rect 69 -21 78 -19
rect 88 -14 97 -12
rect 88 -19 90 -14
rect 95 -19 97 -14
rect 88 -21 97 -19
rect 107 -14 116 -12
rect 107 -19 109 -14
rect 114 -19 116 -14
rect 107 -21 116 -19
rect 126 -14 135 -12
rect 126 -19 128 -14
rect 133 -19 135 -14
rect 126 -21 135 -19
rect 145 -14 154 -12
rect 145 -19 147 -14
rect 152 -19 154 -14
rect 145 -21 154 -19
rect 167 -14 176 -12
rect 167 -19 169 -14
rect 174 -19 176 -14
rect 167 -21 176 -19
rect 191 -14 200 -12
rect 191 -19 193 -14
rect 198 -19 200 -14
rect 191 -21 200 -19
rect 208 -14 217 -12
rect 208 -19 210 -14
rect 215 -19 217 -14
rect 208 -21 217 -19
rect 227 -14 236 -12
rect 227 -19 229 -14
rect 234 -19 236 -14
rect 227 -21 236 -19
rect 246 -14 255 -12
rect 246 -19 248 -14
rect 253 -19 255 -14
rect 246 -21 255 -19
rect 266 -14 275 -12
rect 266 -19 268 -14
rect 273 -19 275 -14
rect 266 -21 275 -19
<< nsubdiff >>
rect -7 102 2 104
rect -7 97 -5 102
rect 0 97 2 102
rect -7 95 2 97
rect 12 102 21 104
rect 12 97 14 102
rect 19 97 21 102
rect 12 95 21 97
rect 31 102 40 104
rect 31 97 33 102
rect 38 97 40 102
rect 31 95 40 97
rect 50 102 59 104
rect 50 97 52 102
rect 57 97 59 102
rect 50 95 59 97
rect 69 102 78 104
rect 69 97 71 102
rect 76 97 78 102
rect 69 95 78 97
rect 91 102 100 104
rect 91 97 93 102
rect 98 97 100 102
rect 91 95 100 97
rect 110 102 119 104
rect 110 97 112 102
rect 117 97 119 102
rect 110 95 119 97
rect 129 102 138 104
rect 129 97 131 102
rect 136 97 138 102
rect 129 95 138 97
rect 148 102 157 104
rect 148 97 150 102
rect 155 97 157 102
rect 148 95 157 97
rect 167 102 176 104
rect 167 97 169 102
rect 174 97 176 102
rect 167 95 176 97
rect 182 102 191 104
rect 182 97 184 102
rect 189 97 191 102
rect 182 95 191 97
rect 199 102 208 104
rect 199 97 201 102
rect 206 97 208 102
rect 199 95 208 97
rect 218 102 227 104
rect 218 97 220 102
rect 225 97 227 102
rect 218 95 227 97
rect 237 102 246 104
rect 237 97 239 102
rect 244 97 246 102
rect 237 95 246 97
rect 256 102 265 104
rect 256 97 258 102
rect 263 97 265 102
rect 256 95 265 97
<< psubdiffcont >>
rect -5 -19 0 -14
rect 14 -19 19 -14
rect 33 -19 38 -14
rect 52 -19 57 -14
rect 71 -19 76 -14
rect 90 -19 95 -14
rect 109 -19 114 -14
rect 128 -19 133 -14
rect 147 -19 152 -14
rect 169 -19 174 -14
rect 193 -19 198 -14
rect 210 -19 215 -14
rect 229 -19 234 -14
rect 248 -19 253 -14
rect 268 -19 273 -14
<< nsubdiffcont >>
rect -5 97 0 102
rect 14 97 19 102
rect 33 97 38 102
rect 52 97 57 102
rect 71 97 76 102
rect 93 97 98 102
rect 112 97 117 102
rect 131 97 136 102
rect 150 97 155 102
rect 169 97 174 102
rect 184 97 189 102
rect 201 97 206 102
rect 220 97 225 102
rect 239 97 244 102
rect 258 97 263 102
<< polysilicon >>
rect 3 86 9 91
rect 45 86 51 91
rect 65 86 71 91
rect 113 86 119 91
rect 142 86 148 91
rect 177 86 183 91
rect 221 86 227 91
rect 250 86 256 91
rect 3 40 9 52
rect 45 50 51 52
rect 38 47 51 50
rect 38 42 40 47
rect 47 42 51 47
rect 38 40 51 42
rect -4 37 9 40
rect -4 32 -2 37
rect 5 32 9 37
rect 65 35 71 52
rect 113 50 119 52
rect -4 30 9 32
rect 3 26 9 30
rect 45 31 71 35
rect 76 48 119 50
rect 76 45 108 48
rect 45 26 51 31
rect 76 26 82 45
rect 106 43 108 45
rect 115 43 119 48
rect 142 44 148 52
rect 106 41 119 43
rect 125 40 148 44
rect 177 42 183 52
rect 221 50 227 52
rect 213 47 227 50
rect 213 45 216 47
rect 125 37 137 40
rect 125 35 130 37
rect 3 21 51 26
rect 3 16 9 21
rect 45 16 51 21
rect 65 21 82 26
rect 113 31 130 35
rect 135 35 137 37
rect 144 35 148 40
rect 135 33 148 35
rect 170 39 183 42
rect 214 42 216 45
rect 223 42 227 47
rect 214 40 227 42
rect 250 39 256 52
rect 170 34 172 39
rect 179 34 183 39
rect 234 36 256 39
rect 233 35 256 36
rect 233 34 238 35
rect 170 32 183 34
rect 65 16 71 21
rect 113 16 119 31
rect 135 25 148 28
rect 135 20 137 25
rect 144 20 148 25
rect 135 18 148 20
rect 142 16 148 18
rect 177 24 183 32
rect 221 32 238 34
rect 221 30 237 32
rect 221 24 227 30
rect 177 19 227 24
rect 243 27 256 30
rect 243 22 245 27
rect 252 22 256 27
rect 243 20 256 22
rect 177 16 183 19
rect 221 16 227 19
rect 250 16 256 20
rect 3 -6 9 -1
rect 45 -6 51 -1
rect 65 -6 71 -1
rect 113 -6 119 -1
rect 142 -6 148 -1
rect 177 -6 183 -1
rect 221 -6 227 -1
rect 250 -6 256 -1
<< polycontact >>
rect 40 42 47 47
rect -2 32 5 37
rect 108 43 115 48
rect 137 35 144 40
rect 216 42 223 47
rect 172 34 179 39
rect 137 20 144 25
rect 245 22 252 27
<< metal1 >>
rect -16 102 283 106
rect -16 97 -5 102
rect 0 97 14 102
rect 19 97 33 102
rect 38 97 52 102
rect 57 97 71 102
rect 76 97 93 102
rect 98 97 112 102
rect 117 97 131 102
rect 136 97 150 102
rect 155 97 169 102
rect 174 97 184 102
rect 189 97 201 102
rect 206 97 220 102
rect 225 97 239 102
rect 244 97 258 102
rect 263 97 283 102
rect -16 92 283 97
rect -5 81 0 92
rect -5 72 0 76
rect 12 81 17 84
rect 12 72 17 76
rect 27 82 39 84
rect 27 81 29 82
rect 27 74 29 76
rect 37 74 39 82
rect 27 72 39 74
rect 52 82 64 84
rect 52 74 54 82
rect 62 74 64 82
rect 52 72 64 74
rect 169 81 174 92
rect 169 72 174 76
rect 186 81 191 84
rect 186 72 191 76
rect 258 83 270 85
rect 258 75 260 83
rect 268 75 270 83
rect 258 73 270 75
rect 73 67 85 69
rect -5 63 0 67
rect -5 55 0 58
rect 12 63 17 67
rect 12 49 17 58
rect 27 63 32 67
rect 12 48 22 49
rect 12 42 14 48
rect 20 42 22 48
rect 12 41 22 42
rect -5 38 5 39
rect -5 32 -3 38
rect 3 37 5 38
rect -5 30 5 32
rect 12 28 17 41
rect 12 27 22 28
rect 12 21 14 27
rect 20 21 22 27
rect -5 9 0 13
rect -5 -7 0 4
rect 12 9 17 21
rect 12 1 17 4
rect 27 9 32 58
rect 56 63 61 67
rect 37 48 51 50
rect 37 42 39 48
rect 46 47 51 48
rect 47 42 51 47
rect 37 39 51 42
rect 27 1 32 4
rect 56 9 61 58
rect 73 59 75 67
rect 83 59 85 67
rect 73 57 85 59
rect 95 67 107 69
rect 95 59 97 67
rect 105 59 107 67
rect 95 57 107 59
rect 122 67 134 69
rect 203 67 215 69
rect 122 59 124 67
rect 132 59 134 67
rect 122 57 134 59
rect 152 63 157 67
rect 56 1 61 4
rect 75 9 80 57
rect 75 1 80 4
rect 95 9 100 57
rect 105 49 119 50
rect 105 43 107 49
rect 113 48 119 49
rect 115 43 119 48
rect 105 42 119 43
rect 95 1 100 4
rect 124 9 129 57
rect 134 41 144 42
rect 134 35 136 41
rect 142 40 144 41
rect 134 33 144 35
rect 134 26 144 27
rect 134 20 136 26
rect 142 25 144 26
rect 134 18 144 20
rect 152 11 157 58
rect 169 63 174 67
rect 169 55 174 58
rect 186 63 191 67
rect 186 49 191 58
rect 203 59 205 67
rect 213 59 215 67
rect 203 57 215 59
rect 231 67 243 69
rect 231 66 233 67
rect 231 61 232 66
rect 231 59 233 61
rect 241 59 243 67
rect 231 57 243 59
rect 186 48 196 49
rect 186 42 188 48
rect 194 42 196 48
rect 186 41 196 42
rect 169 40 179 41
rect 169 34 171 40
rect 177 39 179 40
rect 169 32 179 34
rect 186 27 191 41
rect 186 25 196 27
rect 186 19 188 25
rect 194 19 196 25
rect 124 1 129 4
rect 149 9 160 11
rect 149 2 151 9
rect 158 2 160 9
rect 149 0 160 2
rect 169 9 174 13
rect 169 -7 174 4
rect 186 9 191 19
rect 186 1 191 4
rect 203 9 208 57
rect 213 48 223 49
rect 213 42 215 48
rect 221 47 223 48
rect 213 40 223 42
rect 203 1 208 4
rect 232 9 237 57
rect 242 28 252 29
rect 242 22 244 28
rect 250 27 252 28
rect 242 20 252 22
rect 232 1 237 4
rect 260 9 265 73
rect 260 1 265 4
rect -16 -14 283 -7
rect -16 -19 -5 -14
rect 0 -19 14 -14
rect 19 -19 33 -14
rect 38 -19 52 -14
rect 57 -19 71 -14
rect 76 -19 90 -14
rect 95 -19 109 -14
rect 114 -19 128 -14
rect 133 -19 147 -14
rect 152 -19 169 -14
rect 174 -19 193 -14
rect 198 -19 210 -14
rect 215 -19 229 -14
rect 234 -19 248 -14
rect 253 -19 268 -14
rect 273 -19 283 -14
rect -16 -21 283 -19
<< via1 >>
rect 29 81 37 82
rect 29 76 36 81
rect 36 76 37 81
rect 29 74 37 76
rect 54 81 62 82
rect 54 76 56 81
rect 56 76 61 81
rect 61 76 62 81
rect 54 74 62 76
rect 260 82 268 83
rect 260 77 262 82
rect 262 77 267 82
rect 267 77 268 82
rect 260 75 268 77
rect 14 42 20 48
rect -3 37 3 38
rect -3 32 -2 37
rect -2 32 3 37
rect 14 21 20 27
rect 39 47 46 48
rect 39 42 40 47
rect 40 42 46 47
rect 75 66 83 67
rect 75 61 77 66
rect 77 61 82 66
rect 82 61 83 66
rect 75 59 83 61
rect 97 66 105 67
rect 97 61 99 66
rect 99 61 104 66
rect 104 61 105 66
rect 97 59 105 61
rect 124 59 132 67
rect 107 48 113 49
rect 107 43 108 48
rect 108 43 113 48
rect 136 40 142 41
rect 136 35 137 40
rect 137 35 142 40
rect 136 25 142 26
rect 136 20 137 25
rect 137 20 142 25
rect 205 66 213 67
rect 205 61 207 66
rect 207 61 212 66
rect 212 61 213 66
rect 205 59 213 61
rect 233 66 241 67
rect 233 61 240 66
rect 240 61 241 66
rect 233 59 241 61
rect 188 42 194 48
rect 171 39 177 40
rect 171 34 172 39
rect 172 34 177 39
rect 188 19 194 25
rect 151 2 158 9
rect 215 47 221 48
rect 215 42 216 47
rect 216 42 221 47
rect 244 27 250 28
rect 244 22 245 27
rect 245 22 250 27
<< metal2 >>
rect 27 82 39 84
rect 27 74 29 82
rect 37 74 39 82
rect 27 72 39 74
rect 52 82 64 84
rect 258 83 270 85
rect 258 82 260 83
rect 52 74 54 82
rect 62 75 260 82
rect 268 75 270 83
rect 62 74 64 75
rect 52 72 64 74
rect 258 73 270 75
rect 73 67 85 69
rect 73 59 75 67
rect 83 59 85 67
rect 73 57 85 59
rect 95 67 107 69
rect 95 59 97 67
rect 105 59 107 67
rect 95 57 107 59
rect 122 67 134 69
rect 122 59 124 67
rect 132 63 134 67
rect 203 67 215 69
rect 203 63 205 67
rect 132 59 205 63
rect 213 59 215 67
rect 122 57 215 59
rect 231 67 243 69
rect 231 59 233 67
rect 241 59 243 67
rect 231 57 243 59
rect 37 49 51 50
rect 105 49 119 50
rect 12 48 107 49
rect 12 42 14 48
rect 20 42 39 48
rect 46 43 107 48
rect 113 43 119 49
rect 46 42 119 43
rect 186 48 223 49
rect 186 42 188 48
rect 194 42 215 48
rect 221 42 223 48
rect 12 41 22 42
rect -6 38 5 40
rect 37 39 51 42
rect 134 41 148 42
rect 186 41 223 42
rect -6 32 -3 38
rect 3 32 5 38
rect 134 35 136 41
rect 142 35 148 41
rect 134 33 148 35
rect 168 40 179 41
rect 168 34 171 40
rect 177 34 179 40
rect 168 33 179 34
rect -6 30 5 32
rect 242 28 256 29
rect 12 27 22 28
rect 12 21 14 27
rect 20 26 148 27
rect 20 21 136 26
rect 12 17 22 21
rect 134 20 136 21
rect 142 20 148 26
rect 134 18 148 20
rect 186 25 196 26
rect 242 25 244 28
rect 186 19 188 25
rect 194 22 244 25
rect 250 22 256 28
rect 194 19 256 22
rect 186 17 256 19
rect 149 9 160 11
rect 149 2 151 9
rect 158 2 160 9
rect 149 0 160 2
<< via2 >>
rect -3 32 3 38
rect 136 35 142 41
<< metal3 >>
rect 134 41 148 42
rect -6 39 5 40
rect 134 39 136 41
rect -6 38 136 39
rect -6 32 -3 38
rect 3 35 136 38
rect 142 35 148 41
rect 3 33 148 35
rect 3 32 5 33
rect -6 30 5 32
<< labels >>
rlabel via1 237 63 237 63 3 OUT
port 7 e default output
rlabel via1 102 63 102 63 0 X3
port 4 nsew default input
rlabel via1 79 65 79 65 7 X0
port 3 w default input
rlabel via1 34 79 34 79 7 X1
port 2 w default input
rlabel nsubdiffcont -4 99 -4 99 1 VDD
port 8 n default bidirectional
rlabel psubdiffcont -2 -17 -2 -17 5 VSS
port 9 s default bidirectional
rlabel via1 173 37 173 37 3 C1
port 6 e default input
rlabel via1 154 5 154 5 0 X2
port 5 nsew default input
rlabel via2 -1 34 -1 34 7 C0
port 1 w default input
<< end >>
