* SPICE3 file created from MUX4.ext - technology: gf180mcuC

.option scale=5n

X0 a_1160_210# C1 OUT VDD pfet_03v3 ad=34n pd=0.88m as=23.8n ps=0.48m w=340 l=60
X1 X2 a_250_210# a_590_210# VSS nfet_03v3 ad=22.1n pd=0.6m as=11.9n ps=0.31m w=170 l=60
X2 X0 a_250_210# a_1160_210# VSS nfet_03v3 ad=22.1n pd=0.6m as=12.8n ps=0.33m w=170 l=60
X3 X2 C0 a_590_210# VDD pfet_03v3 ad=44.8n pd=0.96m as=23.8n ps=0.48m w=340 l=60
X4 a_n90_210# C1 VSS VSS nfet_03v3 ad=17n pd=0.54m as=17n ps=0.54m w=170 l=60
X5 X0 C0 a_1160_210# VDD pfet_03v3 ad=44.8n pd=0.96m as=23.8n ps=0.48m w=340 l=60
X6 a_250_210# C0 VSS VSS nfet_03v3 ad=17n pd=0.54m as=17n ps=0.54m w=170 l=60
X7 OUT C1 a_590_210# VSS nfet_03v3 ad=11.9n pd=0.31m as=17n ps=0.54m w=170 l=60
X8 a_n90_210# C1 VDD VDD pfet_03v3 ad=40.8n pd=0.92m as=34n ps=0.88m w=340 l=60
X9 a_250_210# C0 VDD VDD pfet_03v3 ad=34n pd=0.88m as=34n ps=0.88m w=340 l=60
X10 OUT a_n90_210# a_590_210# VDD pfet_03v3 ad=23.8n pd=0.48m as=34.6n ps=0.9m w=340 l=60
X11 a_590_210# C0 X3 VSS nfet_03v3 ad=11.9n pd=0.31m as=17n ps=0.54m w=170 l=60
X12 a_1160_210# C0 X1 VSS nfet_03v3 ad=12.8n pd=0.33m as=17n ps=0.54m w=170 l=60
X13 a_590_210# a_250_210# X3 VDD pfet_03v3 ad=23.8n pd=0.48m as=34.6n ps=0.9m w=340 l=60
X14 a_1160_210# a_n90_210# OUT VSS nfet_03v3 ad=24.1n pd=0.64m as=11.9n ps=0.31m w=170 l=60
X15 a_1160_210# a_250_210# X1 VDD pfet_03v3 ad=23.8n pd=0.48m as=34.6n ps=0.9m w=340 l=60
C0 VDD VSS 5.40677f
