* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__aoi33_1.ext - technology: gf180mcuD

.option scale=5n

X0 a_1310_210# F VSS VSS nfet_03v3 ad=9.35n pd=0.28m as=17n ps=0.54m w=170 l=60
X1 OUT D a_1480_210# VSS nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X2 a_1480_210# E a_1310_210# VSS nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X3 a_1310_720# F OUT VDD pfet_03v3 ad=18.7n pd=0.45m as=34n ps=0.88m w=340 l=60
X4 a_1310_720# D OUT VDD pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X5 a_1820_210# A OUT VSS nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X6 OUT E a_1310_720# VDD pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X7 VSS C a_1990_210# VSS nfet_03v3 ad=17n pd=0.54m as=9.35n ps=0.28m w=170 l=60
X8 a_1990_210# B a_1820_210# VSS nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X9 VDD A a_1310_720# VDD pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X10 VDD C a_1310_720# VDD pfet_03v3 ad=34n pd=0.88m as=18.7n ps=0.45m w=340 l=60
X11 a_1310_720# B VDD VDD pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
C0 a_1310_720# A 0.01969f
C1 OUT F 0.11804f
C2 a_1310_720# B 0.02283f
C3 E OUT 0.05861f
C4 VDD A 0.09996f
C5 VDD B 0.09805f
C6 D a_1310_720# 0.0172f
C7 C B 0.13834f
C8 B a_1990_210# 0.00297f
C9 F A 0
C10 F B 0
C11 VDD D 0.08675f
C12 a_1480_210# D 0.00297f
C13 OUT A 0.1684f
C14 OUT B 0.09467f
C15 F D 0
C16 E D 0.13834f
C17 OUT a_1820_210# 0.00354f
C18 OUT D 0.18649f
C19 A B 0.13834f
C20 VDD a_1310_720# 0.72085f
C21 C a_1310_720# 0.00167f
C22 E a_1310_210# 0.00297f
C23 F a_1310_720# 0.00167f
C24 E a_1310_720# 0.01759f
C25 D A 0.06819f
C26 a_1820_210# A 0.00297f
C27 C VDD 0.10876f
C28 OUT a_1310_210# 0.00232f
C29 VDD F 0.13074f
C30 E VDD 0.08723f
C31 OUT a_1310_720# 0.62324f
C32 C F 0
C33 E F 0.07113f
C34 OUT VDD 0.16592f
C35 OUT a_1480_210# 0.00316f
C36 C OUT 0.10022f
C37 OUT a_1990_210# 0.00297f
C38 OUT VSS 0.42162f
C39 C VSS 0.3984f
C40 B VSS 0.30452f
C41 A VSS 0.30946f
C42 D VSS 0.30954f
C43 E VSS 0.32807f
C44 F VSS 0.39864f
C45 VDD VSS 2.84616f
C46 a_1990_210# VSS 0.00795f **FLOATING
C47 a_1820_210# VSS 0.00738f **FLOATING
C48 a_1480_210# VSS 0.00738f **FLOATING
C49 a_1310_210# VSS 0.00795f **FLOATING
C50 a_1310_720# VSS 0.07075f **FLOATING
