VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__mux4_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__mux4_1 ;
  ORIGIN 0.800 1.050 ;
  SIZE 14.950 BY 6.350 ;
  PIN C0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.295000 ;
    PORT
      LAYER Metal1 ;
        RECT -0.250 1.500 0.250 1.950 ;
        RECT 6.700 1.650 7.200 2.100 ;
      LAYER Metal2 ;
        RECT -0.300 1.500 0.250 2.000 ;
        RECT 6.700 1.650 7.400 2.100 ;
      LAYER Metal3 ;
        RECT -0.300 1.950 0.250 2.000 ;
        RECT 6.700 1.950 7.400 2.100 ;
        RECT -0.300 1.650 7.400 1.950 ;
        RECT -0.300 1.500 0.250 1.650 ;
    END
  END C0
  PIN X1
    DIRECTION INPUT ;
    ANTENNADIFFAREA 2.550000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 3.600 1.950 4.200 ;
        RECT 1.350 0.050 1.600 3.350 ;
      LAYER Metal2 ;
        RECT 1.350 3.600 1.950 4.200 ;
    END
  END X1
  PIN X0
    DIRECTION INPUT ;
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 2.850 4.250 3.450 ;
        RECT 3.750 0.050 4.000 2.850 ;
      LAYER Metal2 ;
        RECT 3.650 2.850 4.250 3.450 ;
    END
  END X0
  PIN X3
    DIRECTION INPUT ;
    ANTENNADIFFAREA 2.550000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 2.850 5.350 3.450 ;
        RECT 4.750 0.050 5.000 2.850 ;
      LAYER Metal2 ;
        RECT 4.750 2.850 5.350 3.450 ;
    END
  END X3
  PIN X2
    DIRECTION INPUT ;
    ANTENNADIFFAREA 1.657500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 0.550 7.850 3.350 ;
        RECT 7.450 0.000 8.000 0.550 ;
      LAYER Metal2 ;
        RECT 7.450 0.000 8.000 0.550 ;
    END
  END X2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 1.600 8.950 2.050 ;
      LAYER Metal2 ;
        RECT 8.400 1.650 8.950 2.050 ;
    END
  END C1
  PIN OUT
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.932500 ;
    PORT
      LAYER Metal1 ;
        RECT 11.550 2.850 12.150 3.450 ;
        RECT 11.600 0.050 11.850 2.850 ;
      LAYER Metal2 ;
        RECT 11.550 2.850 12.150 3.450 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.800 2.100 14.150 4.750 ;
      LAYER Metal1 ;
        RECT -0.800 4.600 14.150 5.300 ;
        RECT -0.250 3.600 0.000 4.600 ;
        RECT 8.450 3.600 8.700 4.600 ;
        RECT -0.250 2.750 0.000 3.350 ;
        RECT 8.450 2.750 8.700 3.350 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT -0.250 -0.350 0.000 0.650 ;
        RECT 8.450 -0.350 8.700 0.650 ;
        RECT -0.800 -1.050 14.150 -0.350 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.600 3.600 0.850 4.200 ;
        RECT 2.600 3.600 3.200 4.200 ;
        RECT 9.300 3.600 9.550 4.200 ;
        RECT 12.900 3.650 13.500 4.250 ;
        RECT 0.600 2.450 0.850 3.350 ;
        RECT 0.600 2.050 1.100 2.450 ;
        RECT 0.600 1.400 0.850 2.050 ;
        RECT 1.850 1.950 2.550 2.500 ;
        RECT 0.600 1.050 1.100 1.400 ;
        RECT 0.600 0.050 0.850 1.050 ;
        RECT 2.800 0.050 3.050 3.350 ;
        RECT 6.100 2.850 6.700 3.450 ;
        RECT 5.250 2.100 5.950 2.500 ;
        RECT 6.200 0.050 6.450 2.850 ;
        RECT 9.300 2.450 9.550 3.350 ;
        RECT 10.150 2.850 10.750 3.450 ;
        RECT 9.300 2.050 9.800 2.450 ;
        RECT 9.300 1.350 9.550 2.050 ;
        RECT 6.700 0.900 7.200 1.350 ;
        RECT 9.300 0.950 9.800 1.350 ;
        RECT 9.300 0.050 9.550 0.950 ;
        RECT 10.150 0.050 10.400 2.850 ;
        RECT 10.650 2.000 11.150 2.450 ;
        RECT 12.100 1.000 12.600 1.450 ;
        RECT 13.000 0.050 13.250 3.650 ;
      LAYER Metal2 ;
        RECT 2.600 4.100 3.200 4.200 ;
        RECT 12.900 4.100 13.500 4.250 ;
        RECT 2.600 3.750 13.500 4.100 ;
        RECT 2.600 3.600 3.200 3.750 ;
        RECT 12.900 3.650 13.500 3.750 ;
        RECT 6.100 3.150 6.700 3.450 ;
        RECT 10.150 3.150 10.750 3.450 ;
        RECT 6.100 2.850 10.750 3.150 ;
        RECT 1.850 2.450 2.550 2.500 ;
        RECT 5.250 2.450 5.950 2.500 ;
        RECT 0.600 2.100 5.950 2.450 ;
        RECT 0.600 2.050 1.100 2.100 ;
        RECT 1.850 1.950 2.550 2.100 ;
        RECT 9.300 2.050 11.150 2.450 ;
        RECT 0.600 1.350 1.100 1.400 ;
        RECT 0.600 1.050 7.400 1.350 ;
        RECT 0.600 0.850 1.100 1.050 ;
        RECT 6.700 0.900 7.400 1.050 ;
        RECT 9.300 1.250 9.800 1.300 ;
        RECT 12.100 1.250 12.800 1.450 ;
        RECT 9.300 0.850 12.800 1.250 ;
  END
END gf180mcu_osu_sc_gp9t3v3__mux4_1
END LIBRARY

