magic
tech gf180mcuD
timestamp 1755575833
<< nwell >>
rect -16 43 283 96
<< nmos >>
rect 3 -4 9 13
rect 45 -4 51 13
rect 65 -4 71 13
rect 113 -4 119 13
rect 142 -4 148 13
rect 177 -4 183 13
rect 221 -4 227 13
rect 250 -4 256 13
<< pmos >>
rect 3 53 9 87
rect 45 53 51 87
rect 65 53 71 87
rect 113 53 119 87
rect 142 53 148 87
rect 177 53 183 87
rect 221 53 227 87
rect 250 53 256 87
<< ndiff >>
rect -7 6 3 13
rect -7 1 -5 6
rect 0 1 3 6
rect -7 -4 3 1
rect 9 6 19 13
rect 9 1 12 6
rect 17 1 19 6
rect 9 -4 19 1
rect 25 6 45 13
rect 25 1 27 6
rect 32 1 45 6
rect 25 -4 45 1
rect 51 6 65 13
rect 51 1 56 6
rect 61 1 65 6
rect 51 -4 65 1
rect 71 6 84 13
rect 71 1 75 6
rect 80 1 84 6
rect 71 -4 84 1
rect 93 6 113 13
rect 93 1 95 6
rect 100 1 113 6
rect 93 -4 113 1
rect 119 6 142 13
rect 119 1 124 6
rect 129 1 142 6
rect 119 -4 142 1
rect 148 6 161 13
rect 148 -1 151 6
rect 158 -1 161 6
rect 148 -4 161 -1
rect 167 6 177 13
rect 167 1 169 6
rect 174 1 177 6
rect 167 -4 177 1
rect 183 6 193 13
rect 183 1 186 6
rect 191 1 193 6
rect 183 -4 193 1
rect 201 6 221 13
rect 201 1 203 6
rect 208 1 221 6
rect 201 -4 221 1
rect 227 6 250 13
rect 227 1 232 6
rect 237 1 250 6
rect 227 -4 250 1
rect 256 6 269 13
rect 256 1 260 6
rect 265 1 269 6
rect 256 -4 269 1
<< pdiff >>
rect -7 82 3 87
rect -7 77 -5 82
rect 0 77 3 82
rect -7 64 3 77
rect -7 59 -5 64
rect 0 59 3 64
rect -7 53 3 59
rect 9 82 19 87
rect 9 77 12 82
rect 17 77 19 82
rect 9 64 19 77
rect 9 59 12 64
rect 17 59 19 64
rect 9 53 19 59
rect 25 82 45 87
rect 25 77 27 82
rect 36 77 45 82
rect 25 64 45 77
rect 25 59 27 64
rect 32 59 45 64
rect 25 53 45 59
rect 51 82 65 87
rect 51 77 56 82
rect 61 77 65 82
rect 51 64 65 77
rect 51 59 56 64
rect 61 59 65 64
rect 51 53 65 59
rect 71 65 87 87
rect 71 60 77 65
rect 82 60 87 65
rect 71 53 87 60
rect 93 65 113 87
rect 93 60 99 65
rect 104 60 113 65
rect 93 53 113 60
rect 119 66 142 87
rect 119 58 124 66
rect 132 58 142 66
rect 119 53 142 58
rect 148 64 161 87
rect 148 59 152 64
rect 157 59 161 64
rect 148 53 161 59
rect 167 82 177 87
rect 167 77 169 82
rect 174 77 177 82
rect 167 64 177 77
rect 167 59 169 64
rect 174 59 177 64
rect 167 53 177 59
rect 183 82 193 87
rect 183 77 186 82
rect 191 77 193 82
rect 183 64 193 77
rect 183 59 186 64
rect 191 59 193 64
rect 183 53 193 59
rect 201 65 221 87
rect 201 60 207 65
rect 212 60 221 65
rect 201 53 221 60
rect 227 63 250 87
rect 227 58 232 63
rect 240 58 250 63
rect 227 53 250 58
rect 256 83 274 87
rect 256 78 262 83
rect 267 78 274 83
rect 256 53 274 78
<< ndiffc >>
rect -5 1 0 6
rect 12 1 17 6
rect 27 1 32 6
rect 56 1 61 6
rect 75 1 80 6
rect 95 1 100 6
rect 124 1 129 6
rect 151 -1 158 6
rect 169 1 174 6
rect 186 1 191 6
rect 203 1 208 6
rect 232 1 237 6
rect 260 1 265 6
<< pdiffc >>
rect -5 77 0 82
rect -5 59 0 64
rect 12 77 17 82
rect 12 59 17 64
rect 27 77 36 82
rect 27 59 32 64
rect 56 77 61 82
rect 56 59 61 64
rect 77 60 82 65
rect 99 60 104 65
rect 124 58 132 66
rect 152 59 157 64
rect 169 77 174 82
rect 169 59 174 64
rect 186 77 191 82
rect 186 59 191 64
rect 207 60 212 65
rect 232 58 240 63
rect 262 78 267 83
<< psubdiff >>
rect -7 -14 2 -12
rect -7 -19 -5 -14
rect 0 -19 2 -14
rect -7 -21 2 -19
rect 12 -14 21 -12
rect 12 -19 14 -14
rect 19 -19 21 -14
rect 12 -21 21 -19
rect 31 -14 40 -12
rect 31 -19 33 -14
rect 38 -19 40 -14
rect 31 -21 40 -19
rect 50 -14 59 -12
rect 50 -19 52 -14
rect 57 -19 59 -14
rect 50 -21 59 -19
rect 69 -14 78 -12
rect 69 -19 71 -14
rect 76 -19 78 -14
rect 69 -21 78 -19
rect 88 -14 97 -12
rect 88 -19 90 -14
rect 95 -19 97 -14
rect 88 -21 97 -19
rect 107 -14 116 -12
rect 107 -19 109 -14
rect 114 -19 116 -14
rect 107 -21 116 -19
rect 126 -14 135 -12
rect 126 -19 128 -14
rect 133 -19 135 -14
rect 126 -21 135 -19
rect 145 -14 154 -12
rect 145 -19 147 -14
rect 152 -19 154 -14
rect 145 -21 154 -19
rect 167 -14 176 -12
rect 167 -19 169 -14
rect 174 -19 176 -14
rect 167 -21 176 -19
rect 191 -14 200 -12
rect 191 -19 193 -14
rect 198 -19 200 -14
rect 191 -21 200 -19
rect 208 -14 217 -12
rect 208 -19 210 -14
rect 215 -19 217 -14
rect 208 -21 217 -19
rect 227 -14 236 -12
rect 227 -19 229 -14
rect 234 -19 236 -14
rect 227 -21 236 -19
rect 246 -14 255 -12
rect 246 -19 248 -14
rect 253 -19 255 -14
rect 246 -21 255 -19
rect 266 -14 275 -12
rect 266 -19 268 -14
rect 273 -19 275 -14
rect 266 -21 275 -19
<< nsubdiff >>
rect -7 103 2 105
rect -7 98 -5 103
rect 0 98 2 103
rect -7 96 2 98
rect 12 103 21 105
rect 12 98 14 103
rect 19 98 21 103
rect 12 96 21 98
rect 31 103 40 105
rect 31 98 33 103
rect 38 98 40 103
rect 31 96 40 98
rect 50 103 59 105
rect 50 98 52 103
rect 57 98 59 103
rect 50 96 59 98
rect 69 103 78 105
rect 69 98 71 103
rect 76 98 78 103
rect 69 96 78 98
rect 91 103 100 105
rect 91 98 93 103
rect 98 98 100 103
rect 91 96 100 98
rect 110 103 119 105
rect 110 98 112 103
rect 117 98 119 103
rect 110 96 119 98
rect 129 103 138 105
rect 129 98 131 103
rect 136 98 138 103
rect 129 96 138 98
rect 148 103 157 105
rect 148 98 150 103
rect 155 98 157 103
rect 148 96 157 98
rect 167 103 176 105
rect 167 98 169 103
rect 174 98 176 103
rect 167 96 176 98
rect 182 103 191 105
rect 182 98 184 103
rect 189 98 191 103
rect 182 96 191 98
rect 199 103 208 105
rect 199 98 201 103
rect 206 98 208 103
rect 199 96 208 98
rect 218 103 227 105
rect 218 98 220 103
rect 225 98 227 103
rect 218 96 227 98
rect 237 103 246 105
rect 237 98 239 103
rect 244 98 246 103
rect 237 96 246 98
rect 256 103 265 105
rect 256 98 258 103
rect 263 98 265 103
rect 256 96 265 98
<< psubdiffcont >>
rect -5 -19 0 -14
rect 14 -19 19 -14
rect 33 -19 38 -14
rect 52 -19 57 -14
rect 71 -19 76 -14
rect 90 -19 95 -14
rect 109 -19 114 -14
rect 128 -19 133 -14
rect 147 -19 152 -14
rect 169 -19 174 -14
rect 193 -19 198 -14
rect 210 -19 215 -14
rect 229 -19 234 -14
rect 248 -19 253 -14
rect 268 -19 273 -14
<< nsubdiffcont >>
rect -5 98 0 103
rect 14 98 19 103
rect 33 98 38 103
rect 52 98 57 103
rect 71 98 76 103
rect 93 98 98 103
rect 112 98 117 103
rect 131 98 136 103
rect 150 98 155 103
rect 169 98 174 103
rect 184 98 189 103
rect 201 98 206 103
rect 220 98 225 103
rect 239 98 244 103
rect 258 98 263 103
<< polysilicon >>
rect 3 87 9 92
rect 45 87 51 92
rect 65 87 71 92
rect 113 87 119 92
rect 142 87 148 92
rect 177 87 183 92
rect 221 87 227 92
rect 250 87 256 92
rect 3 37 9 53
rect 45 51 51 53
rect 38 48 51 51
rect 38 43 40 48
rect 47 43 51 48
rect 38 41 51 43
rect -4 34 9 37
rect -4 29 -2 34
rect 5 29 9 34
rect 65 31 71 53
rect 113 51 119 53
rect -4 27 9 29
rect 3 20 9 27
rect 45 26 71 31
rect 76 48 119 51
rect 76 46 108 48
rect 45 20 51 26
rect 76 20 82 46
rect 106 43 108 46
rect 115 43 119 48
rect 106 41 119 43
rect 142 36 148 53
rect 177 37 183 53
rect 221 51 227 53
rect 213 48 227 51
rect 213 46 216 48
rect 214 43 216 46
rect 223 43 227 48
rect 214 41 227 43
rect 106 33 148 36
rect 106 28 108 33
rect 115 31 148 33
rect 170 34 183 37
rect 250 36 256 53
rect 115 28 119 31
rect 106 26 119 28
rect 170 29 172 34
rect 179 29 183 34
rect 170 27 183 29
rect 3 15 51 20
rect 3 13 9 15
rect 45 13 51 15
rect 65 15 82 20
rect 65 13 71 15
rect 113 13 119 26
rect 135 22 148 25
rect 135 17 137 22
rect 144 17 148 22
rect 135 15 148 17
rect 142 13 148 15
rect 177 20 183 27
rect 221 31 256 36
rect 221 20 227 31
rect 177 15 227 20
rect 243 23 256 26
rect 243 18 245 23
rect 252 18 256 23
rect 243 16 256 18
rect 177 13 183 15
rect 221 13 227 15
rect 250 13 256 16
rect 3 -9 9 -4
rect 45 -9 51 -4
rect 65 -9 71 -4
rect 113 -9 119 -4
rect 142 -9 148 -4
rect 177 -9 183 -4
rect 221 -9 227 -4
rect 250 -9 256 -4
<< polycontact >>
rect 40 43 47 48
rect -2 29 5 34
rect 108 43 115 48
rect 216 43 223 48
rect 108 28 115 33
rect 172 29 179 34
rect 137 17 144 22
rect 245 18 252 23
<< metal1 >>
rect -16 103 283 106
rect -16 98 -5 103
rect 0 98 14 103
rect 19 98 33 103
rect 38 98 52 103
rect 57 98 71 103
rect 76 98 93 103
rect 98 98 112 103
rect 117 98 131 103
rect 136 98 150 103
rect 155 98 169 103
rect 174 98 184 103
rect 189 98 201 103
rect 206 98 220 103
rect 225 98 239 103
rect 244 98 258 103
rect 263 98 283 103
rect -16 94 283 98
rect -5 82 0 94
rect -5 73 0 77
rect 12 82 17 85
rect 12 73 17 77
rect 27 83 39 85
rect 27 82 29 83
rect 27 75 29 77
rect 37 75 39 83
rect 27 73 39 75
rect 52 83 64 85
rect 52 75 54 83
rect 62 75 64 83
rect 52 73 64 75
rect 169 82 174 94
rect 169 73 174 77
rect 186 82 191 85
rect 186 73 191 77
rect 258 84 270 86
rect 258 76 260 84
rect 268 76 270 84
rect 258 74 270 76
rect -5 64 0 68
rect -5 56 0 59
rect 12 64 17 68
rect 12 50 17 59
rect 27 64 32 68
rect 12 49 22 50
rect 12 43 14 49
rect 20 43 22 49
rect 12 42 22 43
rect -5 35 5 36
rect -5 29 -3 35
rect 3 34 5 35
rect -5 27 5 29
rect 12 23 17 42
rect 12 21 22 23
rect 12 15 14 21
rect 20 15 22 21
rect -5 6 0 10
rect -5 -10 0 1
rect 12 6 17 15
rect 12 -2 17 1
rect 27 6 32 59
rect 56 64 61 68
rect 37 49 47 50
rect 37 43 39 49
rect 45 48 47 49
rect 37 41 47 43
rect 27 -2 32 1
rect 56 6 61 59
rect 73 66 85 68
rect 73 58 75 66
rect 83 58 85 66
rect 73 56 85 58
rect 95 66 107 68
rect 95 58 97 66
rect 105 58 107 66
rect 95 56 107 58
rect 122 66 134 68
rect 122 58 124 66
rect 132 58 134 66
rect 122 56 134 58
rect 152 64 157 68
rect 56 -2 61 1
rect 75 6 80 56
rect 75 -2 80 1
rect 95 6 100 56
rect 105 49 115 50
rect 105 43 107 49
rect 113 48 115 49
rect 105 41 115 43
rect 105 34 115 35
rect 105 28 107 34
rect 113 33 115 34
rect 105 26 115 28
rect 95 -2 100 1
rect 124 6 129 56
rect 134 23 144 24
rect 134 17 136 23
rect 142 22 144 23
rect 134 15 144 17
rect 152 8 157 59
rect 169 64 174 68
rect 169 56 174 59
rect 186 64 191 68
rect 186 50 191 59
rect 203 66 215 68
rect 203 58 205 66
rect 213 58 215 66
rect 203 56 215 58
rect 231 64 243 66
rect 231 63 233 64
rect 231 58 232 63
rect 231 56 233 58
rect 241 56 243 64
rect 186 49 196 50
rect 186 43 188 49
rect 194 43 196 49
rect 186 42 196 43
rect 169 35 179 36
rect 169 29 171 35
rect 177 34 179 35
rect 169 27 179 29
rect 186 23 191 42
rect 186 21 196 23
rect 186 15 188 21
rect 194 15 196 21
rect 124 -2 129 1
rect 149 6 160 8
rect 149 -1 151 6
rect 158 -1 160 6
rect 149 -3 160 -1
rect 169 6 174 10
rect 169 -10 174 1
rect 186 6 191 15
rect 186 -2 191 1
rect 203 6 208 56
rect 231 54 243 56
rect 213 49 223 50
rect 213 43 215 49
rect 221 48 223 49
rect 213 41 223 43
rect 203 -2 208 1
rect 232 6 237 54
rect 242 24 252 25
rect 242 18 244 24
rect 250 23 252 24
rect 242 16 252 18
rect 232 -2 237 1
rect 260 6 265 74
rect 260 -2 265 1
rect -16 -14 283 -10
rect -16 -19 -5 -14
rect 0 -19 14 -14
rect 19 -19 33 -14
rect 38 -19 52 -14
rect 57 -19 71 -14
rect 76 -19 90 -14
rect 95 -19 109 -14
rect 114 -19 128 -14
rect 133 -19 147 -14
rect 152 -19 169 -14
rect 174 -19 193 -14
rect 198 -19 210 -14
rect 215 -19 229 -14
rect 234 -19 248 -14
rect 253 -19 268 -14
rect 273 -19 283 -14
rect -16 -21 283 -19
<< via1 >>
rect 29 82 37 83
rect 29 77 36 82
rect 36 77 37 82
rect 29 75 37 77
rect 54 82 62 83
rect 54 77 56 82
rect 56 77 61 82
rect 61 77 62 82
rect 54 75 62 77
rect 260 83 268 84
rect 260 78 262 83
rect 262 78 267 83
rect 267 78 268 83
rect 260 76 268 78
rect 14 43 20 49
rect -3 34 3 35
rect -3 29 -2 34
rect -2 29 3 34
rect 14 15 20 21
rect 39 48 45 49
rect 39 43 40 48
rect 40 43 45 48
rect 75 65 83 66
rect 75 60 77 65
rect 77 60 82 65
rect 82 60 83 65
rect 75 58 83 60
rect 97 65 105 66
rect 97 60 99 65
rect 99 60 104 65
rect 104 60 105 65
rect 97 58 105 60
rect 124 58 132 66
rect 107 48 113 49
rect 107 43 108 48
rect 108 43 113 48
rect 107 33 113 34
rect 107 28 108 33
rect 108 28 113 33
rect 136 22 142 23
rect 136 17 137 22
rect 137 17 142 22
rect 205 65 213 66
rect 205 60 207 65
rect 207 60 212 65
rect 212 60 213 65
rect 205 58 213 60
rect 233 63 241 64
rect 233 58 240 63
rect 240 58 241 63
rect 233 56 241 58
rect 188 43 194 49
rect 171 34 177 35
rect 171 29 172 34
rect 172 29 177 34
rect 188 15 194 21
rect 151 -1 158 6
rect 215 48 221 49
rect 215 43 216 48
rect 216 43 221 48
rect 244 23 250 24
rect 244 18 245 23
rect 245 18 250 23
<< metal2 >>
rect 27 83 39 85
rect 27 75 29 83
rect 37 75 39 83
rect 27 73 39 75
rect 52 83 64 85
rect 258 84 270 86
rect 258 83 260 84
rect 52 75 54 83
rect 62 76 260 83
rect 268 76 270 84
rect 62 75 64 76
rect 52 73 64 75
rect 258 74 270 76
rect 73 66 85 68
rect 73 58 75 66
rect 83 58 85 66
rect 73 56 85 58
rect 95 66 107 68
rect 95 58 97 66
rect 105 58 107 66
rect 95 56 107 58
rect 122 66 134 68
rect 122 58 124 66
rect 132 64 134 66
rect 203 66 215 68
rect 203 64 205 66
rect 132 58 205 64
rect 213 58 215 66
rect 122 56 134 58
rect 203 56 215 58
rect 231 64 243 66
rect 231 56 233 64
rect 241 56 243 64
rect 231 54 243 56
rect 12 49 115 50
rect 12 43 14 49
rect 20 43 39 49
rect 45 43 107 49
rect 113 43 115 49
rect 12 42 115 43
rect 186 49 223 50
rect 186 43 188 49
rect 194 43 215 49
rect 221 43 223 49
rect 186 42 223 43
rect -6 35 5 36
rect 168 35 179 36
rect -6 29 -3 35
rect 3 34 5 35
rect 105 34 119 35
rect 3 29 107 34
rect -6 28 107 29
rect 113 28 119 34
rect 168 29 171 35
rect 177 29 179 35
rect 168 28 179 29
rect 105 27 119 28
rect 242 24 256 25
rect 134 23 148 24
rect 12 21 22 22
rect 12 15 14 21
rect 20 20 22 21
rect 134 20 136 23
rect 20 17 136 20
rect 142 17 148 23
rect 20 15 148 17
rect 12 14 148 15
rect 186 21 196 22
rect 242 21 244 24
rect 186 15 188 21
rect 194 18 244 21
rect 250 18 256 24
rect 194 15 256 18
rect 186 14 256 15
rect 149 6 160 8
rect 149 -1 151 6
rect 158 -1 160 6
rect 149 -3 160 -1
<< labels >>
rlabel nsubdiffcont -4 100 -4 100 1 VDD
rlabel psubdiffcont -2 -17 -2 -17 5 VSS
rlabel via1 0 31 0 31 7 C0
rlabel via1 34 80 34 80 7 X1
rlabel via1 79 64 79 64 7 X0
rlabel via1 102 62 102 62 0 X3
rlabel via1 154 2 154 2 0 X2
rlabel via1 173 32 173 32 3 C1
rlabel via1 237 60 237 60 3 OUT
<< end >>
