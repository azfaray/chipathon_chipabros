magic
tech gf180mcuD
timestamp 1757431385
<< nwell >>
rect 106 63 241 127
<< nmos >>
rect 125 21 131 38
rect 142 21 148 38
rect 159 21 165 38
rect 176 21 182 38
rect 193 21 199 38
rect 210 21 216 38
<< pmos >>
rect 125 72 131 106
rect 142 72 148 106
rect 159 72 165 106
rect 176 72 182 106
rect 193 72 199 106
rect 210 72 216 106
<< ndiff >>
rect 115 36 125 38
rect 115 23 117 36
rect 122 23 125 36
rect 115 21 125 23
rect 131 21 142 38
rect 148 21 159 38
rect 165 36 176 38
rect 165 23 168 36
rect 173 23 176 36
rect 165 21 176 23
rect 182 21 193 38
rect 199 21 210 38
rect 216 36 226 38
rect 216 23 219 36
rect 224 23 226 36
rect 216 21 226 23
<< pdiff >>
rect 115 104 125 106
rect 115 74 117 104
rect 122 74 125 104
rect 115 72 125 74
rect 131 104 142 106
rect 131 85 134 104
rect 139 85 142 104
rect 131 72 142 85
rect 148 94 159 106
rect 148 74 151 94
rect 156 74 159 94
rect 148 72 159 74
rect 165 104 176 106
rect 165 74 168 104
rect 173 74 176 104
rect 165 72 176 74
rect 182 104 193 106
rect 182 84 185 104
rect 190 84 193 104
rect 182 72 193 84
rect 199 104 210 106
rect 199 74 202 104
rect 207 74 210 104
rect 199 72 210 74
rect 216 104 226 106
rect 216 74 219 104
rect 224 74 226 104
rect 216 72 226 74
<< ndiffc >>
rect 117 23 122 36
rect 168 23 173 36
rect 219 23 224 36
<< pdiffc >>
rect 117 74 122 104
rect 134 85 139 104
rect 151 74 156 94
rect 168 74 173 104
rect 185 84 190 104
rect 202 74 207 104
rect 219 74 224 104
<< psubdiff >>
rect 119 12 134 14
rect 119 7 124 12
rect 129 7 134 12
rect 119 5 134 7
rect 143 12 158 14
rect 143 7 148 12
rect 153 7 158 12
rect 143 5 158 7
rect 167 12 182 14
rect 167 7 172 12
rect 177 7 182 12
rect 167 5 182 7
rect 191 12 206 14
rect 191 7 196 12
rect 201 7 206 12
rect 191 5 206 7
rect 215 12 230 14
rect 215 7 220 12
rect 225 7 230 12
rect 215 5 230 7
<< nsubdiff >>
rect 119 120 134 122
rect 119 115 124 120
rect 129 115 134 120
rect 119 113 134 115
rect 143 120 158 122
rect 143 115 148 120
rect 153 115 158 120
rect 143 113 158 115
rect 167 120 182 122
rect 167 115 172 120
rect 177 115 182 120
rect 167 113 182 115
rect 191 120 206 122
rect 191 115 196 120
rect 201 115 206 120
rect 191 113 206 115
rect 215 120 230 122
rect 215 115 220 120
rect 225 115 230 120
rect 215 113 230 115
<< psubdiffcont >>
rect 124 7 129 12
rect 148 7 153 12
rect 172 7 177 12
rect 196 7 201 12
rect 220 7 225 12
<< nsubdiffcont >>
rect 124 115 129 120
rect 148 115 153 120
rect 172 115 177 120
rect 196 115 201 120
rect 220 115 225 120
<< polysilicon >>
rect 125 106 131 111
rect 142 106 148 111
rect 159 106 165 111
rect 176 106 182 111
rect 193 106 199 111
rect 210 106 216 111
rect 125 67 131 72
rect 115 65 131 67
rect 115 59 117 65
rect 123 59 131 65
rect 115 57 131 59
rect 125 38 131 57
rect 142 54 148 72
rect 159 54 165 72
rect 136 52 148 54
rect 136 46 138 52
rect 144 46 148 52
rect 136 44 148 46
rect 153 52 165 54
rect 153 46 155 52
rect 161 46 165 52
rect 153 44 165 46
rect 142 38 148 44
rect 159 38 165 44
rect 176 54 182 72
rect 193 54 199 72
rect 210 54 216 72
rect 176 52 188 54
rect 176 46 180 52
rect 186 46 188 52
rect 176 44 188 46
rect 193 52 205 54
rect 193 46 197 52
rect 203 46 205 52
rect 193 44 205 46
rect 210 52 222 54
rect 210 46 214 52
rect 220 46 222 52
rect 210 44 222 46
rect 176 38 182 44
rect 193 38 199 44
rect 210 38 216 44
rect 125 16 131 21
rect 142 16 148 21
rect 159 16 165 21
rect 176 16 182 21
rect 193 16 199 21
rect 210 16 216 21
<< polycontact >>
rect 117 59 123 65
rect 138 46 144 52
rect 155 46 161 52
rect 180 46 186 52
rect 197 46 203 52
rect 214 46 220 52
<< metal1 >>
rect 106 120 241 127
rect 106 115 124 120
rect 129 115 148 120
rect 153 115 172 120
rect 177 115 196 120
rect 201 115 220 120
rect 225 115 241 120
rect 106 113 241 115
rect 117 104 122 106
rect 134 104 173 106
rect 139 101 168 104
rect 134 83 139 85
rect 151 94 156 96
rect 122 74 151 78
rect 156 74 159 78
rect 117 72 159 74
rect 185 104 190 113
rect 185 82 190 84
rect 202 104 207 106
rect 173 74 202 77
rect 168 72 207 74
rect 219 104 224 113
rect 219 72 224 74
rect 115 59 117 65
rect 123 59 125 65
rect 151 64 156 72
rect 225 64 227 65
rect 151 59 227 64
rect 233 59 235 65
rect 136 46 138 52
rect 144 46 146 52
rect 153 46 155 52
rect 161 46 163 52
rect 117 36 122 38
rect 117 14 122 23
rect 168 36 173 59
rect 178 46 180 52
rect 186 46 188 52
rect 195 46 197 52
rect 203 46 205 52
rect 212 46 214 52
rect 220 46 222 52
rect 168 21 173 23
rect 219 36 224 38
rect 219 14 224 23
rect 106 12 241 14
rect 106 7 124 12
rect 129 7 148 12
rect 153 7 172 12
rect 177 7 196 12
rect 201 7 220 12
rect 225 7 241 12
rect 106 0 241 7
<< via1 >>
rect 117 59 123 65
rect 227 59 233 65
rect 138 46 144 52
rect 155 46 161 52
rect 180 46 186 52
rect 197 46 203 52
rect 214 46 220 52
<< metal2 >>
rect 115 65 125 66
rect 115 59 117 65
rect 123 59 125 65
rect 115 58 125 59
rect 225 65 235 66
rect 225 59 227 65
rect 233 59 235 65
rect 225 58 235 59
rect 136 52 146 53
rect 136 46 138 52
rect 144 46 146 52
rect 136 45 146 46
rect 153 52 163 53
rect 153 46 155 52
rect 161 46 163 52
rect 153 45 163 46
rect 178 52 188 53
rect 178 46 180 52
rect 186 46 188 52
rect 178 45 188 46
rect 195 52 205 53
rect 195 46 197 52
rect 203 46 205 52
rect 195 45 205 46
rect 212 52 222 53
rect 212 46 214 52
rect 220 46 222 52
rect 212 45 222 46
<< labels >>
rlabel nsubdiffcont 124 115 129 120 1 VDD
port 1 n default bidirectional
rlabel metal2 117 59 123 65 7 F
port 5 w default input
rlabel metal2 138 46 144 52 7 E
port 6 w default input
rlabel metal2 155 46 161 52 7 D
port 7 w default input
rlabel metal2 180 46 186 52 7 A
port 4 w default input
rlabel metal2 197 46 203 52 7 B
port 3 w default input
rlabel metal2 214 46 220 52 7 C
port 2 w default input
rlabel psubdiffcont 124 7 129 12 7 VSS
port 9 w default bidirectional
rlabel via1 227 59 233 65 3 OUT
port 8 e default output
<< end >>
