magic
tech gf180mcuD
timestamp 1755780031
use gf180mcu_osu_sc_gp9t3v3__aoi33_1  gf180mcu_osu_sc_gp9t3v3__aoi33_1_0
timestamp 1755277100
transform 1 0 -89 0 1 -50
box 106 0 235 127
use gf180mcu_osu_sc_gp9t3v3__mux4_1  gf180mcu_osu_sc_gp9t3v3__mux4_1_0
timestamp 1755699722
transform 1 0 180 0 1 -50
box -34 0 215 127
use gf180mcu_osu_sc_gp9t3v3__oai33_1  gf180mcu_osu_sc_gp9t3v3__oai33_1_0
timestamp 1755759318
transform 1 0 457 0 1 -47
box -62 -3 67 124
<< end >>
