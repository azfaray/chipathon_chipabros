VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__oai33_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai33_1 ;
  ORIGIN 3.100 0.150 ;
  SIZE 6.450 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -0.450 2.800 0.050 3.100 ;
      LAYER Metal2 ;
        RECT -0.450 2.750 0.050 3.150 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -1.300 2.150 -0.800 2.450 ;
      LAYER Metal2 ;
        RECT -1.300 2.100 -0.800 2.500 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -2.050 2.800 -1.550 3.100 ;
      LAYER Metal2 ;
        RECT -2.050 2.750 -1.550 3.150 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 2.150 0.900 2.450 ;
      LAYER Metal2 ;
        RECT 0.400 2.100 0.900 2.500 ;
    END
  END D
  PIN E
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 2.800 1.750 3.100 ;
      LAYER Metal2 ;
        RECT 1.250 2.750 1.750 3.150 ;
    END
  END E
  PIN F
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 2.150 2.500 2.450 ;
      LAYER Metal2 ;
        RECT 2.000 2.100 2.500 2.500 ;
    END
  END F
  PIN OUT
    ANTENNADIFFAREA 2.592500 ;
    PORT
      LAYER Metal1 ;
        RECT -2.550 3.700 -2.300 5.150 ;
        RECT 2.550 3.700 2.800 5.150 ;
        RECT -2.550 3.450 2.950 3.700 ;
        RECT -2.550 1.900 -2.300 3.450 ;
        RECT 2.700 3.150 2.950 3.450 ;
        RECT 2.650 2.750 3.050 3.150 ;
        RECT -2.550 1.650 -0.600 1.900 ;
        RECT -2.550 0.900 -2.300 1.650 ;
        RECT -0.850 1.300 -0.600 1.650 ;
      LAYER Metal2 ;
        RECT 2.650 2.750 3.050 3.150 ;
    END
  END OUT
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -3.100 3.000 3.350 6.200 ;
      LAYER Metal1 ;
        RECT -3.100 5.500 3.350 6.200 ;
        RECT 0.000 3.950 0.250 5.500 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 0.550 1.100 1.400 ;
        RECT 2.550 0.550 2.800 1.750 ;
        RECT -3.100 -0.150 3.350 0.550 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.000 1.650 1.950 1.900 ;
        RECT -1.700 1.050 -1.450 1.400 ;
        RECT 0.000 1.050 0.250 1.650 ;
        RECT -1.700 0.800 0.250 1.050 ;
        RECT 1.700 0.900 1.950 1.650 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai33_1
END LIBRARY

