* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.ext - technology: gf180mcuD

.option scale=5n

X0 a_510_n10# C1 OUT VDD pfet_03v3 ad=61.2n pd=1.04m as=39.1n ps=0.57m w=340 l=60
X1 X2 C0 a_1190_n10# VDD pfet_03v3 ad=44.2n pd=0.94m as=39.1n ps=0.57m w=340 l=60
X2 a_1190_n10# C0 X3 VSS nfet_03v3 ad=19.55n pd=0.4m as=34n ps=0.74m w=170 l=60
X3 X2 a_90_n10# a_1190_n10# VSS nfet_03v3 ad=22.1n pd=0.6m as=19.55n ps=0.4m w=170 l=60
X4 a_510_n10# a_90_n10# X1 VDD pfet_03v3 ad=23.8n pd=0.48m as=68n ps=1.08m w=340 l=60
X5 OUT C1 a_1190_n10# VSS nfet_03v3 ad=19.55n pd=0.4m as=34n ps=0.74m w=170 l=60
X6 a_510_n10# a_1830_n10# OUT VSS nfet_03v3 ad=22.1n pd=0.6m as=19.55n ps=0.4m w=170 l=60
X7 a_90_n10# C0 VDD VDD pfet_03v3 ad=34n pd=0.88m as=34n ps=0.88m w=340 l=60
X8 a_1830_n10# C1 VSS VSS nfet_03v3 ad=17n pd=0.54m as=17n ps=0.54m w=170 l=60
X9 a_90_n10# C0 VSS VSS nfet_03v3 ad=17n pd=0.54m as=17n ps=0.54m w=170 l=60
X10 a_510_n10# C0 X1 VSS nfet_03v3 ad=11.9n pd=0.31m as=34n ps=0.74m w=170 l=60
X11 X0 C0 a_510_n10# VDD pfet_03v3 ad=54.4n pd=1m as=23.8n ps=0.48m w=340 l=60
X12 OUT a_1830_n10# a_1190_n10# VDD pfet_03v3 ad=39.1n pd=0.57m as=68n ps=1.08m w=340 l=60
X13 a_1190_n10# a_90_n10# X3 VDD pfet_03v3 ad=39.1n pd=0.57m as=68n ps=1.08m w=340 l=60
X14 X0 a_90_n10# a_510_n10# VSS nfet_03v3 ad=22.1n pd=0.6m as=11.9n ps=0.31m w=170 l=60
X15 a_1830_n10# C1 VDD VDD pfet_03v3 ad=34n pd=0.88m as=34n ps=0.88m w=340 l=60
C0 VDD VSS 5.51053f **FLOATING
